-------------------------------------------------------------------------------
-- Title      : Twiddles
-- Project    : 
-------------------------------------------------------------------------------
-- File       : twiddles.vhd
-- Author     : Ola Martin Tiseth Stoevneng  <ola.martin.st@gmail.com>
-- Company    : 
-- Last update: 2014-04-08
-- Platform   : Spartan-6
-------------------------------------------------------------------------------
-- Description: Generated package containing twiddle factors
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author   Description
-- 2014-04-08  1.0      stovneng Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.constants.all;

package twiddles is

  type twat is array(0 to PERDSP*DFT_SIZE-1) of STD_LOGIC_VECTOR(TWLEN-1 downto 0);
  type twa is array(0 to DFT_SIZE/(PERDSP*2)-1) of twat;
  constant TWIDDLES : twa := (
("0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0100000000000000","0100000000000000","0100000000000000",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0010110111010011","0000000011000000","1101001111010011",
"1100000000000000","1101001100101101","0000000001000000","0010110100101101",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","0000000011000000","1100000000000000","0000000001000000",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101",
"0100000000000000","1101001111010011","0000000001000000","0010110111010011",
"1100000000000000","0010110100101101","0000000011000000","1101001100101101"
),
("0100000000000000","0011111111111101","0011111111111010","0011111111110111",
"0011111011110100","0011111011110001","0011110111101110","0011110011101011",
"0011101111101000","0011100111100101","0011100011100010","0011011011100000",
"0011010111011101","0011001111011010","0011000111011000","0010111111010110",
"0010110111010011","0010101011010001","0010100011001111","0010011011001101",
"0010001111001011","0010000011001010","0001111011001000","0001101111000111",
"0001100011000101","0001010111000100","0001001011000011","0000111111000010",
"0000110011000010","0000100111000001","0000011011000001","0000001111000001",
"0000000011000000","1111110111000001","1111101011000001","1111011111000001",
"1111010011000010","1111000111000010","1110111011000011","1110101111000100",
"1110100011000101","1110010111000111","1110001011001000","1110000011001010",
"1101110111001011","1101101011001101","1101100011001111","1101011011010001",
"1101001111010011","1101000111010110","1100111111011000","1100110111011010",
"1100101111011101","1100101011100000","1100100011100010","1100011111100101",
"1100010111101000","1100010011101011","1100001111101110","1100001011110001",
"1100001011110100","1100000111110111","1100000111111010","1100000111111101",
"1100000000000000","1100000100000011","1100000100000110","1100000100001001",
"1100001000001100","1100001000001111","1100001100010010","1100010000010101",
"1100010100011000","1100011100011011","1100100000011110","1100101000100000",
"1100101100100011","1100110100100110","1100111100101000","1101000100101010",
"1101001100101101","1101011000101111","1101100000110001","1101101000110011",
"1101110100110101","1110000000110110","1110001000111000","1110010100111001",
"1110100000111011","1110101100111100","1110111000111101","1111000100111110",
"1111010000111110","1111011100111111","1111101000111111","1111110100111111",
"0000000001000000","0000001100111111","0000011000111111","0000100100111111",
"0000110000111110","0000111100111110","0001001000111101","0001010100111100",
"0001100000111011","0001101100111001","0001111000111000","0010000000110110",
"0010001100110101","0010011000110011","0010100000110001","0010101000101111",
"0010110100101101","0010111100101010","0011000100101000","0011001100100110",
"0011010100100011","0011011000100000","0011100000011110","0011100100011011",
"0011101100011000","0011110000010101","0011110100010010","0011111000001111",
"0011111000001100","0011111100001001","0011111100000110","0011111100000011",
"0100000000000000","0010101011010001","1111101011000001","1100110111011010",
"1100001000001100","1110000000110110","0001001000111101","0011100100011011",
"0011101111101000","0001010111000100","1110001011001000","1100001011110001",
"1100101100100011","1111011100111111","0010100000110001","0011111100000011",
"0010110111010011","1111110111000001","1100111111011000","1100000100001001",
"1101110100110101","0000111100111110","0011100000011110","0011110011101011",
"0001100011000101","1110010111000111","1100001111101110","1100101000100000",
"1111010000111110","0010011000110011","0011111100000110","0010111111010110",
"0000000011000000","1101000111010110","1100000100000110","1101101000110011",
"0000110000111110","0011011000100000","0011110111101110","0001101111000111",
"1110100011000101","1100010011101011","1100100000011110","1111000100111110",
"0010001100110101","0011111100001001","0011000111011000","0000001111000001",
"1101001111010011","1100000100000011","1101100000110001","0000100100111111",
"0011010100100011","0011111011110001","0001111011001000","1110101111000100",
"1100010111101000","1100011100011011","1110111000111101","0010000000110110",
"0011111000001100","0011001111011010","0000011011000001","1101011011010001",
"1100000000000000","1101011000101111","0000011000111111","0011001100100110",
"0011111011110100","0010000011001010","1110111011000011","1100011111100101",
"1100010100011000","1110101100111100","0001111000111000","0011111000001111",
"0011010111011101","0000100111000001","1101100011001111","1100000111111101",
"1101001100101101","0000001100111111","0011000100101000","0011111111110111",
"0010001111001011","1111000111000010","1100100011100010","1100010000010101",
"1110100000111011","0001101100111001","0011110100010010","0011011011100000",
"0000110011000010","1101101011001101","1100000111111010","1101000100101010",
"0000000001000000","0010111100101010","0011111111111010","0010011011001101",
"1111010011000010","1100101011100000","1100001100010010","1110010100111001",
"0001100000111011","0011110000010101","0011100011100010","0000111111000010",
"1101110111001011","1100000111110111","1100111100101000","1111110100111111",
"0010110100101101","0011111111111101","0010100011001111","1111011111000001",
"1100101111011101","1100001000001111","1110001000111000","0001010100111100",
"0011101100011000","0011100111100101","0001001011000011","1110000011001010",
"1100001011110100","1100110100100110","1111101000111111","0010101000101111",
"0100000000000000","1111110111000001","1100000100000110","0000100100111111",
"0011111011110100","1111000111000010","1100001100010010","0001010100111100",
"0011101111101000","1110010111000111","1100100000011110","0010000000110110",
"0011010111011101","1101101011001101","1100111100101000","0010101000101111",
"0010110111010011","1101000111010110","1101100000110001","0011001100100110",
"0010001111001011","1100101011100000","1110001000111000","0011100100011011",
"0001100011000101","1100010011101011","1110111000111101","0011111000001111",
"0000110011000010","1100000111110111","1111101000111111","0011111100000011",
"0000000011000000","1100000100000011","0000011000111111","0011111111110111",
"1111010011000010","1100001000001111","0001001000111101","0011110011101011",
"1110100011000101","1100011100011011","0001111000111000","0011011011100000",
"1101110111001011","1100110100100110","0010100000110001","0010111111010110",
"1101001111010011","1101011000101111","0011000100101000","0010011011001101",
"1100101111011101","1110000000110110","0011100000011110","0001101111000111",
"1100010111101000","1110101100111100","0011110100010010","0000111111000010",
"1100001011110100","1111011100111111","0011111100000110","0000001111000001",
"1100000000000000","0000001100111111","0011111111111010","1111011111000001",
"1100001000001100","0000111100111110","0011110111101110","1110101111000100",
"1100010100011000","0001101100111001","0011100011100010","1110000011001010",
"1100101100100011","0010011000110011","0011000111011000","1101011011010001",
"1101001100101101","0010111100101010","0010100011001111","1100110111011010",
"1101110100110101","0011011000100000","0001111011001000","1100011111100101",
"1110100000111011","0011110000010101","0001001011000011","1100001011110001",
"1111010000111110","0011111100001001","0000011011000001","1100000111111101",
"0000000001000000","0011111111111101","1111101011000001","1100000100001001",
"0000110000111110","0011111011110001","1110111011000011","1100010000010101",
"0001100000111011","0011100111100101","1110001011001000","1100101000100000",
"0010001100110101","0011001111011010","1101100011001111","1101000100101010",
"0010110100101101","0010101011010001","1100111111011000","1101101000110011",
"0011010100100011","0010000011001010","1100100011100010","1110010100111001",
"0011101100011000","0001010111000100","1100001111101110","1111000100111110",
"0011111000001100","0000100111000001","1100000111111010","1111110100111111",
"0100000000000000","1101000111010110","0000011000111111","0010011011001101",
"1100001000001100","0011011000100000","1110111011000011","1110010100111001",
"0011101111101000","1100010011101011","0001111000111000","0000111111000010",
"1100101100100011","0011111100001001","1101100011001111","1111110100111111",
"0010110111010011","1100000100000011","0011000100101000","1111011111000001",
"1101110100110101","0011111011110001","1100100011100010","0001010100111100",
"0001100011000101","1100011100011011","0011110100010010","1110000011001010",
"1111010000111110","0011001111011010","1100000111111010","0010101000101111",
"0000000011000000","1101011000101111","0011111111111010","1100110111011010",
"0000110000111110","0010000011001010","1100001100010010","0011100100011011",
"1110100011000101","1110101100111100","0011100011100010","1100001011110001",
"0010001100110101","0000100111000001","1100111100101000","0011111100000011",
"1101001111010011","0000001100111111","0010100011001111","1100000100001001",
"0011010100100011","1111000111000010","1110001000111000","0011110011101011",
"1100010111101000","0001101100111001","0001001011000011","1100101000100000",
"0011111000001100","1101101011001101","1111101000111111","0010111111010110",
"1100000000000000","0010111100101010","1111101011000001","1101101000110011",
"0011111011110100","1100101011100000","0001001000111101","0001101111000111",
"1100010100011000","0011110000010101","1110001011001000","1111000100111110",
"0011010111011101","1100000111110111","0010100000110001","0000001111000001",
"1101001100101101","0011111111111101","1100111111011000","0000100100111111",
"0010001111001011","1100001000001111","0011100000011110","1110101111000100",
"1110100000111011","0011100111100101","1100001111101110","0010000000110110",
"0000110011000010","1100110100100110","0011111100000110","1101011011010001",
"0000000001000000","0010101011010001","1100000100000110","0011001100100110",
"1111010011000010","1110000000110110","0011110111101110","1100011111100101",
"0001100000111011","0001010111000100","1100100000011110","0011111000001111",
"1101110111001011","1111011100111111","0011000111011000","1100000111111101",
"0010110100101101","1111110111000001","1101100000110001","0011111111110111",
"1100101111011101","0000111100111110","0001111011001000","1100010000010101",
"0011101100011000","1110010111000111","1110111000111101","0011011011100000",
"1100001011110100","0010011000110011","0000011011000001","1101000100101010"
),
("0100000000000000","0011111111111010","0011111011110100","0011110111101110",
"0011101111101000","0011100011100010","0011010111011101","0011000111011000",
"0010110111010011","0010100011001111","0010001111001011","0001111011001000",
"0001100011000101","0001001011000011","0000110011000010","0000011011000001",
"0000000011000000","1111101011000001","1111010011000010","1110111011000011",
"1110100011000101","1110001011001000","1101110111001011","1101100011001111",
"1101001111010011","1100111111011000","1100101111011101","1100100011100010",
"1100010111101000","1100001111101110","1100001011110100","1100000111111010",
"1100000000000000","1100000100000110","1100001000001100","1100001100010010",
"1100010100011000","1100100000011110","1100101100100011","1100111100101000",
"1101001100101101","1101100000110001","1101110100110101","1110001000111000",
"1110100000111011","1110111000111101","1111010000111110","1111101000111111",
"0000000001000000","0000011000111111","0000110000111110","0001001000111101",
"0001100000111011","0001111000111000","0010001100110101","0010100000110001",
"0010110100101101","0011000100101000","0011010100100011","0011100000011110",
"0011101100011000","0011110100010010","0011111000001100","0011111100000110",
"0100000000000000","0011111111111010","0011111011110100","0011110111101110",
"0011101111101000","0011100011100010","0011010111011101","0011000111011000",
"0010110111010011","0010100011001111","0010001111001011","0001111011001000",
"0001100011000101","0001001011000011","0000110011000010","0000011011000001",
"0000000011000000","1111101011000001","1111010011000010","1110111011000011",
"1110100011000101","1110001011001000","1101110111001011","1101100011001111",
"1101001111010011","1100111111011000","1100101111011101","1100100011100010",
"1100010111101000","1100001111101110","1100001011110100","1100000111111010",
"1100000000000000","1100000100000110","1100001000001100","1100001100010010",
"1100010100011000","1100100000011110","1100101100100011","1100111100101000",
"1101001100101101","1101100000110001","1101110100110101","1110001000111000",
"1110100000111011","1110111000111101","1111010000111110","1111101000111111",
"0000000001000000","0000011000111111","0000110000111110","0001001000111101",
"0001100000111011","0001111000111000","0010001100110101","0010100000110001",
"0010110100101101","0011000100101000","0011010100100011","0011100000011110",
"0011101100011000","0011110100010010","0011111000001100","0011111100000110",
"0100000000000000","0010100011001111","1111010011000010","1100100011100010",
"1100010100011000","1110111000111101","0010001100110101","0011111100000110",
"0010110111010011","1111101011000001","1100101111011101","1100001100010010",
"1110100000111011","0001111000111000","0011111000001100","0011000111011000",
"0000000011000000","1100111111011000","1100001000001100","1110001000111000",
"0001100000111011","0011110100010010","0011010111011101","0000011011000001",
"1101001111010011","1100000100000110","1101110100110101","0001001000111101",
"0011101100011000","0011100011100010","0000110011000010","1101100011001111",
"1100000000000000","1101100000110001","0000110000111110","0011100000011110",
"0011101111101000","0001001011000011","1101110111001011","1100000111111010",
"1101001100101101","0000011000111111","0011010100100011","0011110111101110",
"0001100011000101","1110001011001000","1100001011110100","1100111100101000",
"0000000001000000","0011000100101000","0011111011110100","0001111011001000",
"1110100011000101","1100001111101110","1100101100100011","1111101000111111",
"0010110100101101","0011111111111010","0010001111001011","1110111011000011",
"1100010111101000","1100100000011110","1111010000111110","0010100000110001",
"0100000000000000","0010100011001111","1111010011000010","1100100011100010",
"1100010100011000","1110111000111101","0010001100110101","0011111100000110",
"0010110111010011","1111101011000001","1100101111011101","1100001100010010",
"1110100000111011","0001111000111000","0011111000001100","0011000111011000",
"0000000011000000","1100111111011000","1100001000001100","1110001000111000",
"0001100000111011","0011110100010010","0011010111011101","0000011011000001",
"1101001111010011","1100000100000110","1101110100110101","0001001000111101",
"0011101100011000","0011100011100010","0000110011000010","1101100011001111",
"1100000000000000","1101100000110001","0000110000111110","0011100000011110",
"0011101111101000","0001001011000011","1101110111001011","1100000111111010",
"1101001100101101","0000011000111111","0011010100100011","0011110111101110",
"0001100011000101","1110001011001000","1100001011110100","1100111100101000",
"0000000001000000","0011000100101000","0011111011110100","0001111011001000",
"1110100011000101","1100001111101110","1100101100100011","1111101000111111",
"0010110100101101","0011111111111010","0010001111001011","1110111011000011",
"1100010111101000","1100100000011110","1111010000111110","0010100000110001",
"0100000000000000","1111101011000001","1100001000001100","0001001000111101",
"0011101111101000","1110001011001000","1100101100100011","0010100000110001",
"0010110111010011","1100111111011000","1101110100110101","0011100000011110",
"0001100011000101","1100001111101110","1111010000111110","0011111100000110",
"0000000011000000","1100000100000110","0000110000111110","0011110111101110",
"1110100011000101","1100100000011110","0010001100110101","0011000111011000",
"1101001111010011","1101100000110001","0011010100100011","0001111011001000",
"1100010111101000","1110111000111101","0011111000001100","0000011011000001",
"1100000000000000","0000011000111111","0011111011110100","1110111011000011",
"1100010100011000","0001111000111000","0011010111011101","1101100011001111",
"1101001100101101","0011000100101000","0010001111001011","1100100011100010",
"1110100000111011","0011110100010010","0000110011000010","1100000111111010",
"0000000001000000","0011111111111010","1111010011000010","1100001100010010",
"0001100000111011","0011100011100010","1101110111001011","1100111100101000",
"0010110100101101","0010100011001111","1100101111011101","1110001000111000",
"0011101100011000","0001001011000011","1100001011110100","1111101000111111",
"0100000000000000","1111101011000001","1100001000001100","0001001000111101",
"0011101111101000","1110001011001000","1100101100100011","0010100000110001",
"0010110111010011","1100111111011000","1101110100110101","0011100000011110",
"0001100011000101","1100001111101110","1111010000111110","0011111100000110",
"0000000011000000","1100000100000110","0000110000111110","0011110111101110",
"1110100011000101","1100100000011110","0010001100110101","0011000111011000",
"1101001111010011","1101100000110001","0011010100100011","0001111011001000",
"1100010111101000","1110111000111101","0011111000001100","0000011011000001",
"1100000000000000","0000011000111111","0011111011110100","1110111011000011",
"1100010100011000","0001111000111000","0011010111011101","1101100011001111",
"1101001100101101","0011000100101000","0010001111001011","1100100011100010",
"1110100000111011","0011110100010010","0000110011000010","1100000111111010",
"0000000001000000","0011111111111010","1111010011000010","1100001100010010",
"0001100000111011","0011100011100010","1101110111001011","1100111100101000",
"0010110100101101","0010100011001111","1100101111011101","1110001000111000",
"0011101100011000","0001001011000011","1100001011110100","1111101000111111",
"0100000000000000","1100111111011000","0000110000111110","0001111011001000",
"1100010100011000","0011110100010010","1101110111001011","1111101000111111",
"0010110111010011","1100000100000110","0011010100100011","1110111011000011",
"1110100000111011","0011100011100010","1100001011110100","0010100000110001",
"0000000011000000","1101100000110001","0011111011110100","1100100011100010",
"0001100000111011","0001001011000011","1100101100100011","0011111100000110",
"1101001111010011","0000011000111111","0010001111001011","1100001100010010",
"0011101100011000","1110001011001000","1111010000111110","0011000111011000",
"1100000000000000","0011000100101000","1111010011000010","1110001000111000",
"0011101111101000","1100001111101110","0010001100110101","0000011011000001",
"1101001100101101","0011111111111010","1100101111011101","0001001000111101",
"0001100011000101","1100100000011110","0011111000001100","1101100011001111",
"0000000001000000","0010100011001111","1100001000001100","0011100000011110",
"1110100011000101","1110111000111101","0011010111011101","1100000111111010",
"0010110100101101","1111101011000001","1101110100110101","0011110111101110",
"1100010111101000","0001111000111000","0000110011000010","1100111100101000",
"0100000000000000","1100111111011000","0000110000111110","0001111011001000",
"1100010100011000","0011110100010010","1101110111001011","1111101000111111",
"0010110111010011","1100000100000110","0011010100100011","1110111011000011",
"1110100000111011","0011100011100010","1100001011110100","0010100000110001",
"0000000011000000","1101100000110001","0011111011110100","1100100011100010",
"0001100000111011","0001001011000011","1100101100100011","0011111100000110",
"1101001111010011","0000011000111111","0010001111001011","1100001100010010",
"0011101100011000","1110001011001000","1111010000111110","0011000111011000",
"1100000000000000","0011000100101000","1111010011000010","1110001000111000",
"0011101111101000","1100001111101110","0010001100110101","0000011011000001",
"1101001100101101","0011111111111010","1100101111011101","0001001000111101",
"0001100011000101","1100100000011110","0011111000001100","1101100011001111",
"0000000001000000","0010100011001111","1100001000001100","0011100000011110",
"1110100011000101","1110111000111101","0011010111011101","1100000111111010",
"0010110100101101","1111101011000001","1101110100110101","0011110111101110",
"1100010111101000","0001111000111000","0000110011000010","1100111100101000"
),
("0100000000000000","0011111111110111","0011110111101110","0011100111100101",
"0011010111011101","0010111111010110","0010100011001111","0010000011001010",
"0001100011000101","0000111111000010","0000011011000001","1111110111000001",
"1111010011000010","1110101111000100","1110001011001000","1101101011001101",
"1101001111010011","1100110111011010","1100100011100010","1100010011101011",
"1100001011110100","1100000111111101","1100000100000110","1100001000001111",
"1100010100011000","1100101000100000","1100111100101000","1101011000101111",
"1101110100110101","1110010100111001","1110111000111101","1111011100111111",
"0000000001000000","0000100100111111","0001001000111101","0001101100111001",
"0010001100110101","0010101000101111","0011000100101000","0011011000100000",
"0011101100011000","0011111000001111","0011111100000110","0011111111111101",
"0011111011110100","0011110011101011","0011100011100010","0011001111011010",
"0010110111010011","0010011011001101","0001111011001000","0001010111000100",
"0000110011000010","0000001111000001","1111101011000001","1111000111000010",
"1110100011000101","1110000011001010","1101100011001111","1101000111010110",
"1100101111011101","1100011111100101","1100001111101110","1100000111110111",
"1100000000000000","1100000100001001","1100001100010010","1100011100011011",
"1100101100100011","1101000100101010","1101100000110001","1110000000110110",
"1110100000111011","1111000100111110","1111101000111111","0000001100111111",
"0000110000111110","0001010100111100","0001111000111000","0010011000110011",
"0010110100101101","0011001100100110","0011100000011110","0011110000010101",
"0011111000001100","0011111100000011","0011111111111010","0011111011110001",
"0011101111101000","0011011011100000","0011000111011000","0010101011010001",
"0010001111001011","0001101111000111","0001001011000011","0000100111000001",
"0000000011000000","1111011111000001","1110111011000011","1110010111000111",
"1101110111001011","1101011011010001","1100111111011000","1100101011100000",
"1100010111101000","1100001011110001","1100000111111010","1100000100000011",
"1100001000001100","1100010000010101","1100100000011110","1100110100100110",
"1101001100101101","1101101000110011","1110001000111000","1110101100111100",
"1111010000111110","1111110100111111","0000011000111111","0000111100111110",
"0001100000111011","0010000000110110","0010100000110001","0010111100101010",
"0011010100100011","0011100100011011","0011110100010010","0011111100001001",
"0100000000000000","0010011011001101","1110111011000011","1100010011101011",
"1100101100100011","1111110100111111","0011000100101000","0011111011110001",
"0001100011000101","1110000011001010","1100000111111010","1101011000101111",
"0000110000111110","0011100100011011","0011100011100010","0000100111000001",
"1101001111010011","1100000100001001","1110001000111000","0001101100111001",
"0011111000001100","0010111111010110","1111101011000001","1100101011100000",
"1100010100011000","1111000100111110","0010100000110001","0011111111111101",
"0010001111001011","1110101111000100","1100001111101110","1100110100100110",
"0000000001000000","0011001100100110","0011110111101110","0001010111000100",
"1101110111001011","1100000111111101","1101100000110001","0000111100111110",
"0011101100011000","0011011011100000","0000011011000001","1101000111010110",
"1100001000001100","1110010100111001","0001111000111000","0011111100001001",
"0010110111010011","1111011111000001","1100100011100010","1100011100011011",
"1111010000111110","0010101000101111","0011111111111010","0010000011001010",
"1110100011000101","1100001011110001","1100111100101000","0000001100111111",
"0011010100100011","0011110011101011","0001001011000011","1101101011001101",
"1100000000000000","1101101000110011","0001001000111101","0011110000010101",
"0011010111011101","0000001111000001","1100111111011000","1100001000001111",
"1110100000111011","0010000000110110","0011111100000110","0010101011010001",
"1111010011000010","1100011111100101","1100100000011110","1111011100111111",
"0010110100101101","0011111111110111","0001111011001000","1110010111000111",
"1100001011110100","1101000100101010","0000011000111111","0011011000100000",
"0011101111101000","0000111111000010","1101100011001111","1100000100000011",
"1101110100110101","0001010100111100","0011110100010010","0011001111011010",
"0000000011000000","1100110111011010","1100001100010010","1110101100111100",
"0010001100110101","0011111100000011","0010100011001111","1111000111000010",
"1100010111101000","1100101000100000","1111101000111111","0010111100101010",
"0011111011110100","0001101111000111","1110001011001000","1100000111110111",
"1101001100101101","0000100100111111","0011100000011110","0011100111100101",
"0000110011000010","1101011011010001","1100000100000110","1110000000110110",
"0001100000111011","0011111000001111","0011000111011000","1111110111000001",
"1100101111011101","1100010000010101","1110111000111101","0010011000110011",
"0100000000000000","1111011111000001","1100001100010010","0001101100111001",
"0011010111011101","1101011011010001","1101100000110001","0011011000100000",
"0001100011000101","1100001011110001","1111101000111111","0011111111111101",
"1111010011000010","1100010000010101","0001111000111000","0011001111011010",
"1101001111010011","1101101000110011","0011100000011110","0001010111000100",
"1100001011110100","1111110100111111","0011111111111010","1111000111000010",
"1100010100011000","0010000000110110","0011000111011000","1101000111010110",
"1101110100110101","0011100100011011","0001001011000011","1100000111110111",
"0000000001000000","0011111111110111","1110111011000011","1100011100011011",
"0010001100110101","0010111111010110","1100111111011000","1110000000110110",
"0011101100011000","0000111111000010","1100000111111010","0000001100111111",
"0011111011110100","1110101111000100","1100100000011110","0010011000110011",
"0010110111010011","1100110111011010","1110001000111000","0011110000010101",
"0000110011000010","1100000111111101","0000011000111111","0011111011110001",
"1110100011000101","1100101000100000","0010100000110001","0010101011010001",
"1100101111011101","1110010100111001","0011110100010010","0000100111000001",
"1100000000000000","0000100100111111","0011110111101110","1110010111000111",
"1100101100100011","0010101000101111","0010100011001111","1100101011100000",
"1110100000111011","0011111000001111","0000011011000001","1100000100000011",
"0000110000111110","0011110011101011","1110001011001000","1100110100100110",
"0010110100101101","0010011011001101","1100100011100010","1110101100111100",
"0011111000001100","0000001111000001","1100000100000110","0000111100111110",
"0011101111101000","1110000011001010","1100111100101000","0010111100101010",
"0010001111001011","1100011111100101","1110111000111101","0011111100001001",
"0000000011000000","1100000100001001","0001001000111101","0011100111100101",
"1101110111001011","1101000100101010","0011000100101000","0010000011001010",
"1100010111101000","1111000100111110","0011111100000110","1111110111000001",
"1100001000001100","0001010100111100","0011100011100010","1101101011001101",
"1101001100101101","0011001100100110","0001111011001000","1100010011101011",
"1111010000111110","0011111100000011","1111101011000001","1100001000001111",
"0001100000111011","0011011011100000","1101100011001111","1101011000101111",
"0011010100100011","0001101111000111","1100001111101110","1111011100111111",
"0100000000000000","1100110111011010","0001001000111101","0001010111000100",
"1100101100100011","0011111100000011","1100111111011000","0000111100111110",
"0001100011000101","1100101000100000","0011111100000110","1101000111010110",
"0000110000111110","0001101111000111","1100100000011110","0011111100001001",
"1101001111010011","0000100100111111","0001111011001000","1100011100011011",
"0011111000001100","1101011011010001","0000011000111111","0010000011001010",
"1100010100011000","0011111000001111","1101100011001111","0000001100111111",
"0010001111001011","1100010000010101","0011110100010010","1101101011001101",
"0000000001000000","0010011011001101","1100001100010010","0011110000010101",
"1101110111001011","1111110100111111","0010100011001111","1100001000001111",
"0011101100011000","1110000011001010","1111101000111111","0010101011010001",
"1100001000001100","0011100100011011","1110001011001000","1111011100111111",
"0010110111010011","1100000100001001","0011100000011110","1110010111000111",
"1111010000111110","0010111111010110","1100000100000110","0011011000100000",
"1110100011000101","1111000100111110","0011000111011000","1100000100000011",
"0011010100100011","1110101111000100","1110111000111101","0011001111011010",
"1100000000000000","0011001100100110","1110111011000011","1110101100111100",
"0011010111011101","1100000111111101","0011000100101000","1111000111000010",
"1110100000111011","0011011011100000","1100000111111010","0010111100101010",
"1111010011000010","1110010100111001","0011100011100010","1100000111110111",
"0010110100101101","1111011111000001","1110001000111000","0011100111100101",
"1100001011110100","0010101000101111","1111101011000001","1110000000110110",
"0011101111101000","1100001011110001","0010100000110001","1111110111000001",
"1101110100110101","0011110011101011","1100001111101110","0010011000110011",
"0000000011000000","1101101000110011","0011110111101110","1100010011101011",
"0010001100110101","0000001111000001","1101100000110001","0011111011110001",
"1100010111101000","0010000000110110","0000011011000001","1101011000101111",
"0011111011110100","1100011111100101","0001111000111000","0000100111000001",
"1101001100101101","0011111111110111","1100100011100010","0001101100111001",
"0000110011000010","1101000100101010","0011111111111010","1100101011100000",
"0001100000111011","0000111111000010","1100111100101000","0011111111111101",
"1100101111011101","0001010100111100","0001001011000011","1100110100100110"
),
("0100000000000000","0011111011110100","0011101111101000","0011010111011101",
"0010110111010011","0010001111001011","0001100011000101","0000110011000010",
"0000000011000000","1111010011000010","1110100011000101","1101110111001011",
"1101001111010011","1100101111011101","1100010111101000","1100001011110100",
"1100000000000000","1100001000001100","1100010100011000","1100101100100011",
"1101001100101101","1101110100110101","1110100000111011","1111010000111110",
"0000000001000000","0000110000111110","0001100000111011","0010001100110101",
"0010110100101101","0011010100100011","0011101100011000","0011111000001100",
"0100000000000000","0011111011110100","0011101111101000","0011010111011101",
"0010110111010011","0010001111001011","0001100011000101","0000110011000010",
"0000000011000000","1111010011000010","1110100011000101","1101110111001011",
"1101001111010011","1100101111011101","1100010111101000","1100001011110100",
"1100000000000000","1100001000001100","1100010100011000","1100101100100011",
"1101001100101101","1101110100110101","1110100000111011","1111010000111110",
"0000000001000000","0000110000111110","0001100000111011","0010001100110101",
"0010110100101101","0011010100100011","0011101100011000","0011111000001100",
"0100000000000000","0011111011110100","0011101111101000","0011010111011101",
"0010110111010011","0010001111001011","0001100011000101","0000110011000010",
"0000000011000000","1111010011000010","1110100011000101","1101110111001011",
"1101001111010011","1100101111011101","1100010111101000","1100001011110100",
"1100000000000000","1100001000001100","1100010100011000","1100101100100011",
"1101001100101101","1101110100110101","1110100000111011","1111010000111110",
"0000000001000000","0000110000111110","0001100000111011","0010001100110101",
"0010110100101101","0011010100100011","0011101100011000","0011111000001100",
"0100000000000000","0011111011110100","0011101111101000","0011010111011101",
"0010110111010011","0010001111001011","0001100011000101","0000110011000010",
"0000000011000000","1111010011000010","1110100011000101","1101110111001011",
"1101001111010011","1100101111011101","1100010111101000","1100001011110100",
"1100000000000000","1100001000001100","1100010100011000","1100101100100011",
"1101001100101101","1101110100110101","1110100000111011","1111010000111110",
"0000000001000000","0000110000111110","0001100000111011","0010001100110101",
"0010110100101101","0011010100100011","0011101100011000","0011111000001100",
"0100000000000000","0010001111001011","1110100011000101","1100001011110100",
"1101001100101101","0000110000111110","0011101100011000","0011010111011101",
"0000000011000000","1100101111011101","1100010100011000","1111010000111110",
"0010110100101101","0011111011110100","0001100011000101","1101110111001011",
"1100000000000000","1101110100110101","0001100000111011","0011111000001100",
"0010110111010011","1111010011000010","1100010111101000","1100101100100011",
"0000000001000000","0011010100100011","0011101111101000","0000110011000010",
"1101001111010011","1100001000001100","1110100000111011","0010001100110101",
"0100000000000000","0010001111001011","1110100011000101","1100001011110100",
"1101001100101101","0000110000111110","0011101100011000","0011010111011101",
"0000000011000000","1100101111011101","1100010100011000","1111010000111110",
"0010110100101101","0011111011110100","0001100011000101","1101110111001011",
"1100000000000000","1101110100110101","0001100000111011","0011111000001100",
"0010110111010011","1111010011000010","1100010111101000","1100101100100011",
"0000000001000000","0011010100100011","0011101111101000","0000110011000010",
"1101001111010011","1100001000001100","1110100000111011","0010001100110101",
"0100000000000000","0010001111001011","1110100011000101","1100001011110100",
"1101001100101101","0000110000111110","0011101100011000","0011010111011101",
"0000000011000000","1100101111011101","1100010100011000","1111010000111110",
"0010110100101101","0011111011110100","0001100011000101","1101110111001011",
"1100000000000000","1101110100110101","0001100000111011","0011111000001100",
"0010110111010011","1111010011000010","1100010111101000","1100101100100011",
"0000000001000000","0011010100100011","0011101111101000","0000110011000010",
"1101001111010011","1100001000001100","1110100000111011","0010001100110101",
"0100000000000000","0010001111001011","1110100011000101","1100001011110100",
"1101001100101101","0000110000111110","0011101100011000","0011010111011101",
"0000000011000000","1100101111011101","1100010100011000","1111010000111110",
"0010110100101101","0011111011110100","0001100011000101","1101110111001011",
"1100000000000000","1101110100110101","0001100000111011","0011111000001100",
"0010110111010011","1111010011000010","1100010111101000","1100101100100011",
"0000000001000000","0011010100100011","0011101111101000","0000110011000010",
"1101001111010011","1100001000001100","1110100000111011","0010001100110101",
"0100000000000000","1111010011000010","1100010100011000","0010001100110101",
"0010110111010011","1100101111011101","1110100000111011","0011111000001100",
"0000000011000000","1100001000001100","0001100000111011","0011010111011101",
"1101001111010011","1101110100110101","0011101100011000","0000110011000010",
"1100000000000000","0000110000111110","0011101111101000","1101110111001011",
"1101001100101101","0011010100100011","0001100011000101","1100001011110100",
"0000000001000000","0011111011110100","1110100011000101","1100101100100011",
"0010110100101101","0010001111001011","1100010111101000","1111010000111110",
"0100000000000000","1111010011000010","1100010100011000","0010001100110101",
"0010110111010011","1100101111011101","1110100000111011","0011111000001100",
"0000000011000000","1100001000001100","0001100000111011","0011010111011101",
"1101001111010011","1101110100110101","0011101100011000","0000110011000010",
"1100000000000000","0000110000111110","0011101111101000","1101110111001011",
"1101001100101101","0011010100100011","0001100011000101","1100001011110100",
"0000000001000000","0011111011110100","1110100011000101","1100101100100011",
"0010110100101101","0010001111001011","1100010111101000","1111010000111110",
"0100000000000000","1111010011000010","1100010100011000","0010001100110101",
"0010110111010011","1100101111011101","1110100000111011","0011111000001100",
"0000000011000000","1100001000001100","0001100000111011","0011010111011101",
"1101001111010011","1101110100110101","0011101100011000","0000110011000010",
"1100000000000000","0000110000111110","0011101111101000","1101110111001011",
"1101001100101101","0011010100100011","0001100011000101","1100001011110100",
"0000000001000000","0011111011110100","1110100011000101","1100101100100011",
"0010110100101101","0010001111001011","1100010111101000","1111010000111110",
"0100000000000000","1111010011000010","1100010100011000","0010001100110101",
"0010110111010011","1100101111011101","1110100000111011","0011111000001100",
"0000000011000000","1100001000001100","0001100000111011","0011010111011101",
"1101001111010011","1101110100110101","0011101100011000","0000110011000010",
"1100000000000000","0000110000111110","0011101111101000","1101110111001011",
"1101001100101101","0011010100100011","0001100011000101","1100001011110100",
"0000000001000000","0011111011110100","1110100011000101","1100101100100011",
"0010110100101101","0010001111001011","1100010111101000","1111010000111110",
"0100000000000000","1100101111011101","0001100000111011","0000110011000010",
"1101001100101101","0011111011110100","1100010111101000","0010001100110101",
"0000000011000000","1101110100110101","0011101111101000","1100001011110100",
"0010110100101101","1111010011000010","1110100000111011","0011010111011101",
"1100000000000000","0011010100100011","1110100011000101","1111010000111110",
"0010110111010011","1100001000001100","0011101100011000","1101110111001011",
"0000000001000000","0010001111001011","1100010100011000","0011111000001100",
"1101001111010011","0000110000111110","0001100011000101","1100101100100011",
"0100000000000000","1100101111011101","0001100000111011","0000110011000010",
"1101001100101101","0011111011110100","1100010111101000","0010001100110101",
"0000000011000000","1101110100110101","0011101111101000","1100001011110100",
"0010110100101101","1111010011000010","1110100000111011","0011010111011101",
"1100000000000000","0011010100100011","1110100011000101","1111010000111110",
"0010110111010011","1100001000001100","0011101100011000","1101110111001011",
"0000000001000000","0010001111001011","1100010100011000","0011111000001100",
"1101001111010011","0000110000111110","0001100011000101","1100101100100011",
"0100000000000000","1100101111011101","0001100000111011","0000110011000010",
"1101001100101101","0011111011110100","1100010111101000","0010001100110101",
"0000000011000000","1101110100110101","0011101111101000","1100001011110100",
"0010110100101101","1111010011000010","1110100000111011","0011010111011101",
"1100000000000000","0011010100100011","1110100011000101","1111010000111110",
"0010110111010011","1100001000001100","0011101100011000","1101110111001011",
"0000000001000000","0010001111001011","1100010100011000","0011111000001100",
"1101001111010011","0000110000111110","0001100011000101","1100101100100011",
"0100000000000000","1100101111011101","0001100000111011","0000110011000010",
"1101001100101101","0011111011110100","1100010111101000","0010001100110101",
"0000000011000000","1101110100110101","0011101111101000","1100001011110100",
"0010110100101101","1111010011000010","1110100000111011","0011010111011101",
"1100000000000000","0011010100100011","1110100011000101","1111010000111110",
"0010110111010011","1100001000001100","0011101100011000","1101110111001011",
"0000000001000000","0010001111001011","1100010100011000","0011111000001100",
"1101001111010011","0000110000111110","0001100011000101","1100101100100011"
),
("0100000000000000","0011111011110001","0011100011100010","0010111111010110",
"0010001111001011","0001010111000100","0000011011000001","1111011111000001",
"1110100011000101","1101101011001101","1100111111011000","1100011111100101",
"1100001011110100","1100000100000011","1100001100010010","1100101000100000",
"1101001100101101","1110000000110110","1110111000111101","1111110100111111",
"0000110000111110","0001101100111001","0010100000110001","0011001100100110",
"0011101100011000","0011111100001001","0011111111111010","0011110011101011",
"0011010111011101","0010101011010001","0001111011001000","0000111111000010",
"0000000011000000","1111000111000010","1110001011001000","1101011011010001",
"1100101111011101","1100010011101011","1100000111111010","1100000100001001",
"1100010100011000","1100110100100110","1101100000110001","1110010100111001",
"1111010000111110","0000001100111111","0001001000111101","0010000000110110",
"0010110100101101","0011011000100000","0011110100010010","0011111100000011",
"0011111011110100","0011100111100101","0011000111011000","0010011011001101",
"0001100011000101","0000100111000001","1111101011000001","1110101111000100",
"1101110111001011","1101000111010110","1100100011100010","1100001011110001",
"1100000000000000","1100001000001111","1100100000011110","1101000100101010",
"1101110100110101","1110101100111100","1111101000111111","0000100100111111",
"0001100000111011","0010011000110011","0011000100101000","0011100100011011",
"0011111000001100","0011111111111101","0011110111101110","0011011011100000",
"0010110111010011","0010000011001010","0001001011000011","0000001111000001",
"1111010011000010","1110010111000111","1101100011001111","1100110111011010",
"1100010111101000","1100000111110111","1100000100000110","1100010000010101",
"1100101100100011","1101011000101111","1110001000111000","1111000100111110",
"0000000001000000","0000111100111110","0001111000111000","0010101000101111",
"0011010100100011","0011110000010101","0011111100000110","0011111111110111",
"0011101111101000","0011001111011010","0010100011001111","0001101111000111",
"0000110011000010","1111110111000001","1110111011000011","1110000011001010",
"1101001111010011","1100101011100000","1100001111101110","1100000111111101",
"1100001000001100","1100011100011011","1100111100101000","1101101000110011",
"1110100000111011","1111011100111111","0000011000111111","0001010100111100",
"0010001100110101","0010111100101010","0011100000011110","0011111000001111",
"0100000000000000","0010000011001010","1110001011001000","1100000111111101",
"1101110100110101","0001101100111001","0011111100000110","0010011011001101",
"1110100011000101","1100000111110111","1101100000110001","0001010100111100",
"0011111000001100","0010101011010001","1110111011000011","1100001011110001",
"1101001100101101","0000111100111110","0011110100010010","0010111111010110",
"1111010011000010","1100010011101011","1100111100101000","0000100100111111",
"0011101100011000","0011001111011010","1111101011000001","1100011111100101",
"1100101100100011","0000001100111111","0011100000011110","0011011011100000",
"0000000011000000","1100101011100000","1100100000011110","1111110100111111",
"0011010100100011","0011100111100101","0000011011000001","1100110111011010",
"1100010100011000","1111011100111111","0011000100101000","0011110011101011",
"0000110011000010","1101000111010110","1100001100010010","1111000100111110",
"0010110100101101","0011111011110001","0001001011000011","1101011011010001",
"1100001000001100","1110101100111100","0010100000110001","0011111111110111",
"0001100011000101","1101101011001101","1100000100000110","1110010100111001",
"0010001100110101","0011111111111101","0001111011001000","1110000011001010",
"1100000000000000","1110000000110110","0001111000111000","0011111100000011",
"0010001111001011","1110010111000111","1100000111111010","1101101000110011",
"0001100000111011","0011111100001001","0010100011001111","1110101111000100",
"1100001011110100","1101011000101111","0001001000111101","0011111000001111",
"0010110111010011","1111000111000010","1100001111101110","1101000100101010",
"0000110000111110","0011110000010101","0011000111011000","1111011111000001",
"1100010111101000","1100110100100110","0000011000111111","0011100100011011",
"0011010111011101","1111110111000001","1100100011100010","1100101000100000",
"0000000001000000","0011011000100000","0011100011100010","0000001111000001",
"1100101111011101","1100011100011011","1111101000111111","0011001100100110",
"0011101111101000","0000100111000001","1100111111011000","1100010000010101",
"1111010000111110","0010111100101010","0011110111101110","0000111111000010",
"1101001111010011","1100001000001111","1110111000111101","0010101000101111",
"0011111011110100","0001010111000100","1101100011001111","1100000100001001",
"1110100000111011","0010011000110011","0011111111111010","0001101111000111",
"1101110111001011","1100000100000011","1110001000111000","0010000000110110",
"0100000000000000","1111000111000010","1100100000011110","0010101000101111",
"0010001111001011","1100010011101011","1111101000111111","0011111111110111",
"1110100011000101","1100110100100110","0011000100101000","0001101111000111",
"1100001011110100","0000001100111111","0011110111101110","1110000011001010",
"1101001100101101","0011011000100000","0001001011000011","1100000111111101",
"0000110000111110","0011100111100101","1101100011001111","1101101000110011",
"0011101100011000","0000100111000001","1100000100000110","0001010100111100",
"0011010111011101","1101000111010110","1110001000111000","0011111000001111",
"0000000011000000","1100001000001111","0001111000111000","0010111111010110",
"1100101111011101","1110101100111100","0011111100000110","1111011111000001",
"1100010100011000","0010011000110011","0010100011001111","1100011111100101",
"1111010000111110","0011111111111101","1110111011000011","1100101000100000",
"0010110100101101","0010000011001010","1100001111101110","1111110100111111",
"0011111011110100","1110010111000111","1100111100101000","0011001100100110",
"0001100011000101","1100000111110111","0000011000111111","0011110011101011",
"1101110111001011","1101011000101111","0011100000011110","0000111111000010",
"1100000000000000","0000111100111110","0011100011100010","1101011011010001",
"1101110100110101","0011110000010101","0000011011000001","1100000100001001",
"0001100000111011","0011001111011010","1100111111011000","1110010100111001",
"0011111000001100","1111110111000001","1100001100010010","0010000000110110",
"0010110111010011","1100101011100000","1110111000111101","0011111100000011",
"1111010011000010","1100011100011011","0010100000110001","0010011011001101",
"1100010111101000","1111011100111111","0011111111111010","1110101111000100",
"1100101100100011","0010111100101010","0001111011001000","1100001011110001",
"0000000001000000","0011111011110001","1110001011001000","1101000100101010",
"0011010100100011","0001010111000100","1100000111111010","0000100100111111",
"0011101111101000","1101101011001101","1101100000110001","0011100100011011",
"0000110011000010","1100000100000011","0001001000111101","0011011011100000",
"1101001111010011","1110000000110110","0011110100010010","0000001111000001",
"1100001000001100","0001101100111001","0011000111011000","1100110111011010",
"1110100000111011","0011111100001001","1111101011000001","1100010000010101",
"0010001100110101","0010101011010001","1100100011100010","1111000100111110",
"0100000000000000","1100101011100000","0001111000111000","0000001111000001",
"1101110100110101","0011100111100101","1100000111111010","0011001100100110",
"1110100011000101","1111011100111111","0010100011001111","1100010000010101",
"0011111000001100","1101000111010110","0001001000111101","0000111111000010",
"1101001100101101","0011111011110001","1100001111101110","0010101000101111",
"1111010011000010","1110101100111100","0011000111011000","1100000100001001",
"0011101100011000","1101101011001101","0000011000111111","0001101111000111",
"1100101100100011","0011111111111101","1100100011100010","0010000000110110",
"0000000011000000","1110000000110110","0011100011100010","1100000111111101",
"0011010100100011","1110010111000111","1111101000111111","0010011011001101",
"1100010100011000","0011111100001001","1100111111011000","0001010100111100",
"0000110011000010","1101011000101111","0011110111101110","1100001011110001",
"0010110100101101","1111000111000010","1110111000111101","0010111111010110",
"1100001000001100","0011110000010101","1101100011001111","0000100100111111",
"0001100011000101","1100110100100110","0011111111111010","1100011111100101",
"0010001100110101","1111110111000001","1110001000111000","0011011011100000",
"1100000000000000","0011011000100000","1110001011001000","1111110100111111",
"0010001111001011","1100011100011011","0011111100000110","1100110111011010",
"0001100000111011","0000100111000001","1101100000110001","0011110011101011",
"1100001011110100","0010111100101010","1110111011000011","1111000100111110",
"0010110111010011","1100001000001111","0011110100010010","1101011011010001",
"0000110000111110","0001010111000100","1100111100101000","0011111111110111",
"1100010111101000","0010011000110011","1111101011000001","1110010100111001",
"0011010111011101","1100000100000011","0011100000011110","1110000011001010",
"0000000001000000","0010000011001010","1100100000011110","0011111100000011",
"1100101111011101","0001101100111001","0000011011000001","1101101000110011",
"0011101111101000","1100000111110111","0011000100101000","1110101111000100",
"1111010000111110","0010101011010001","1100001100010010","0011111000001111",
"1101001111010011","0000111100111110","0001001011000011","1101000100101010",
"0011111011110100","1100010011101011","0010100000110001","1111011111000001",
"1110100000111011","0011001111011010","1100000100000110","0011100100011011",
"1101110111001011","0000001100111111","0001111011001000","1100101000100000"
),
("0100000000000000","0011110111101110","0011010111011101","0010100011001111",
"0001100011000101","0000011011000001","1111010011000010","1110001011001000",
"1101001111010011","1100100011100010","1100001011110100","1100000100000110",
"1100010100011000","1100111100101000","1101110100110101","1110111000111101",
"0000000001000000","0001001000111101","0010001100110101","0011000100101000",
"0011101100011000","0011111100000110","0011111011110100","0011100011100010",
"0010110111010011","0001111011001000","0000110011000010","1111101011000001",
"1110100011000101","1101100011001111","1100101111011101","1100001111101110",
"1100000000000000","1100001100010010","1100101100100011","1101100000110001",
"1110100000111011","1111101000111111","0000110000111110","0001111000111000",
"0010110100101101","0011100000011110","0011111000001100","0011111111111010",
"0011101111101000","0011000111011000","0010001111001011","0001001011000011",
"0000000011000000","1110111011000011","1101110111001011","1100111111011000",
"1100010111101000","1100000111111010","1100001000001100","1100100000011110",
"1101001100101101","1110001000111000","1111010000111110","0000011000111111",
"0001100000111011","0010100000110001","0011010100100011","0011110100010010",
"0100000000000000","0011110111101110","0011010111011101","0010100011001111",
"0001100011000101","0000011011000001","1111010011000010","1110001011001000",
"1101001111010011","1100100011100010","1100001011110100","1100000100000110",
"1100010100011000","1100111100101000","1101110100110101","1110111000111101",
"0000000001000000","0001001000111101","0010001100110101","0011000100101000",
"0011101100011000","0011111100000110","0011111011110100","0011100011100010",
"0010110111010011","0001111011001000","0000110011000010","1111101011000001",
"1110100011000101","1101100011001111","1100101111011101","1100001111101110",
"1100000000000000","1100001100010010","1100101100100011","1101100000110001",
"1110100000111011","1111101000111111","0000110000111110","0001111000111000",
"0010110100101101","0011100000011110","0011111000001100","0011111111111010",
"0011101111101000","0011000111011000","0010001111001011","0001001011000011",
"0000000011000000","1110111011000011","1101110111001011","1100111111011000",
"1100010111101000","1100000111111010","1100001000001100","1100100000011110",
"1101001100101101","1110001000111000","1111010000111110","0000011000111111",
"0001100000111011","0010100000110001","0011010100100011","0011110100010010",
"0100000000000000","0001111011001000","1101110111001011","1100000100000110",
"1110100000111011","0010100000110001","0011111011110100","0001001011000011",
"1101001111010011","1100001100010010","1111010000111110","0011000100101000",
"0011101111101000","0000011011000001","1100101111011101","1100100000011110",
"0000000001000000","0011100000011110","0011010111011101","1111101011000001",
"1100010111101000","1100111100101000","0000110000111110","0011110100010010",
"0010110111010011","1110111011000011","1100001011110100","1101100000110001",
"0001100000111011","0011111100000110","0010001111001011","1110001011001000",
"1100000000000000","1110001000111000","0010001100110101","0011111111111010",
"0001100011000101","1101100011001111","1100001000001100","1110111000111101",
"0010110100101101","0011110111101110","0000110011000010","1100111111011000",
"1100010100011000","1111101000111111","0011010100100011","0011100011100010",
"0000000011000000","1100100011100010","1100101100100011","0000011000111111",
"0011101100011000","0011000111011000","1111010011000010","1100001111101110",
"1101001100101101","0001001000111101","0011111000001100","0010100011001111",
"1110100011000101","1100000111111010","1101110100110101","0001111000111000",
"0100000000000000","0001111011001000","1101110111001011","1100000100000110",
"1110100000111011","0010100000110001","0011111011110100","0001001011000011",
"1101001111010011","1100001100010010","1111010000111110","0011000100101000",
"0011101111101000","0000011011000001","1100101111011101","1100100000011110",
"0000000001000000","0011100000011110","0011010111011101","1111101011000001",
"1100010111101000","1100111100101000","0000110000111110","0011110100010010",
"0010110111010011","1110111011000011","1100001011110100","1101100000110001",
"0001100000111011","0011111100000110","0010001111001011","1110001011001000",
"1100000000000000","1110001000111000","0010001100110101","0011111111111010",
"0001100011000101","1101100011001111","1100001000001100","1110111000111101",
"0010110100101101","0011110111101110","0000110011000010","1100111111011000",
"1100010100011000","1111101000111111","0011010100100011","0011100011100010",
"0000000011000000","1100100011100010","1100101100100011","0000011000111111",
"0011101100011000","0011000111011000","1111010011000010","1100001111101110",
"1101001100101101","0001001000111101","0011111000001100","0010100011001111",
"1110100011000101","1100000111111010","1101110100110101","0001111000111000",
"0100000000000000","1110111011000011","1100101100100011","0011000100101000",
"0001100011000101","1100000111111010","0000110000111110","0011100011100010",
"1101001111010011","1110001000111000","0011111000001100","1111101011000001",
"1100010100011000","0010100000110001","0010001111001011","1100001111101110",
"0000000001000000","0011110111101110","1101110111001011","1101100000110001",
"0011101100011000","0000011011000001","1100001000001100","0001111000111000",
"0010110111010011","1100100011100010","1111010000111110","0011111111111010",
"1110100011000101","1100111100101000","0011010100100011","0001001011000011",
"1100000000000000","0001001000111101","0011010111011101","1100111111011000",
"1110100000111011","0011111100000110","1111010011000010","1100100000011110",
"0010110100101101","0001111011001000","1100001011110100","0000011000111111",
"0011101111101000","1101100011001111","1101110100110101","0011110100010010",
"0000000011000000","1100001100010010","0010001100110101","0010100011001111",
"1100010111101000","1111101000111111","0011111011110100","1110001011001000",
"1101001100101101","0011100000011110","0000110011000010","1100000100000110",
"0001100000111011","0011000111011000","1100101111011101","1110111000111101",
"0100000000000000","1110111011000011","1100101100100011","0011000100101000",
"0001100011000101","1100000111111010","0000110000111110","0011100011100010",
"1101001111010011","1110001000111000","0011111000001100","1111101011000001",
"1100010100011000","0010100000110001","0010001111001011","1100001111101110",
"0000000001000000","0011110111101110","1101110111001011","1101100000110001",
"0011101100011000","0000011011000001","1100001000001100","0001111000111000",
"0010110111010011","1100100011100010","1111010000111110","0011111111111010",
"1110100011000101","1100111100101000","0011010100100011","0001001011000011",
"1100000000000000","0001001000111101","0011010111011101","1100111111011000",
"1110100000111011","0011111100000110","1111010011000010","1100100000011110",
"0010110100101101","0001111011001000","1100001011110100","0000011000111111",
"0011101111101000","1101100011001111","1101110100110101","0011110100010010",
"0000000011000000","1100001100010010","0010001100110101","0010100011001111",
"1100010111101000","1111101000111111","0011111011110100","1110001011001000",
"1101001100101101","0011100000011110","0000110011000010","1100000100000110",
"0001100000111011","0011000111011000","1100101111011101","1110111000111101",
"0100000000000000","1100100011100010","0010001100110101","1111101011000001",
"1110100000111011","0011000111011000","1100001000001100","0011110100010010",
"1101001111010011","0001001000111101","0000110011000010","1101100000110001",
"0011101111101000","1100000111111010","0011010100100011","1110001011001000",
"0000000001000000","0001111011001000","1100101100100011","0011111111111010",
"1100010111101000","0010100000110001","1111010011000010","1110111000111101",
"0010110111010011","1100001100010010","0011111000001100","1100111111011000",
"0001100000111011","0000011011000001","1101110100110101","0011100011100010",
"1100000000000000","0011100000011110","1101110111001011","0000011000111111",
"0001100011000101","1100111100101000","0011111011110100","1100001111101110",
"0010110100101101","1110111011000011","1111010000111110","0010100011001111",
"1100010100011000","0011111100000110","1100101111011101","0001111000111000",
"0000000011000000","1110001000111000","0011010111011101","1100000100000110",
"0011101100011000","1101100011001111","0000110000111110","0001001011000011",
"1101001100101101","0011110111101110","1100001011110100","0011000100101000",
"1110100011000101","1111101000111111","0010001111001011","1100100000011110",
"0100000000000000","1100100011100010","0010001100110101","1111101011000001",
"1110100000111011","0011000111011000","1100001000001100","0011110100010010",
"1101001111010011","0001001000111101","0000110011000010","1101100000110001",
"0011101111101000","1100000111111010","0011010100100011","1110001011001000",
"0000000001000000","0001111011001000","1100101100100011","0011111111111010",
"1100010111101000","0010100000110001","1111010011000010","1110111000111101",
"0010110111010011","1100001100010010","0011111000001100","1100111111011000",
"0001100000111011","0000011011000001","1101110100110101","0011100011100010",
"1100000000000000","0011100000011110","1101110111001011","0000011000111111",
"0001100011000101","1100111100101000","0011111011110100","1100001111101110",
"0010110100101101","1110111011000011","1111010000111110","0010100011001111",
"1100010100011000","0011111100000110","1100101111011101","0001111000111000",
"0000000011000000","1110001000111000","0011010111011101","1100000100000110",
"0011101100011000","1101100011001111","0000110000111110","0001001011000011",
"1101001100101101","0011110111101110","1100001011110100","0011000100101000",
"1110100011000101","1111101000111111","0010001111001011","1100100000011110"
),
("0100000000000000","0011110011101011","0011000111011000","0010000011001010",
"0000110011000010","1111011111000001","1110001011001000","1101000111010110",
"1100010111101000","1100000111111101","1100001100010010","1100110100100110",
"1101110100110101","1111000100111110","0000011000111111","0001101100111001",
"0010110100101101","0011100100011011","0011111100000110","0011111011110001",
"0011010111011101","0010011011001101","0001001011000011","1111110111000001",
"1110100011000101","1101011011010001","1100100011100010","1100000111110111",
"1100001000001100","1100101000100000","1101100000110001","1110101100111100",
"0000000001000000","0001010100111100","0010100000110001","0011011000100000",
"0011111000001100","0011111111110111","0011100011100010","0010101011010001",
"0001100011000101","0000001111000001","1110111011000011","1101101011001101",
"1100101111011101","1100001011110001","1100000100000110","1100011100011011",
"1101001100101101","1110010100111001","1111101000111111","0000111100111110",
"0010001100110101","0011001100100110","0011110100010010","0011111111111101",
"0011101111101000","0010111111010110","0001111011001000","0000100111000001",
"1111010011000010","1110000011001010","1100111111011000","1100010011101011",
"1100000000000000","1100010000010101","1100111100101000","1110000000110110",
"1111010000111110","0000100100111111","0001111000111000","0010111100101010",
"0011101100011000","0011111100000011","0011110111101110","0011001111011010",
"0010001111001011","0000111111000010","1111101011000001","1110010111000111",
"1101001111010011","1100011111100101","1100000111111010","1100001000001111",
"1100101100100011","1101101000110011","1110111000111101","0000001100111111",
"0001100000111011","0010101000101111","0011100000011110","0011111100001001",
"0011111011110100","0011011011100000","0010100011001111","0001010111000100",
"0000000011000000","1110101111000100","1101100011001111","1100101011100000",
"1100001011110100","1100000100001001","1100100000011110","1101011000101111",
"1110100000111011","1111110100111111","0001001000111101","0010011000110011",
"0011010100100011","0011111000001111","0011111111111010","0011100111100101",
"0010110111010011","0001101111000111","0000011011000001","1111000111000010",
"1101110111001011","1100110111011010","1100001111101110","1100000100000011",
"1100010100011000","1101000100101010","1110001000111000","1111011100111111",
"0000110000111110","0010000000110110","0011000100101000","0011110000010101",
"0100000000000000","0001101111000111","1101100011001111","1100001000001111",
"1111010000111110","0011001100100110","0011100011100010","1111110111000001",
"1100010111101000","1101000100101010","0001001000111101","0011111100001001",
"0010001111001011","1110000011001010","1100000100000110","1110101100111100",
"0010110100101101","0011110011101011","0000011011000001","1100101011100000",
"1100101100100011","0000100100111111","0011110100010010","0010101011010001",
"1110100011000101","1100000111111101","1110001000111000","0010011000110011",
"0011111011110100","0000111111000010","1100111111011000","1100011100011011",
"0000000001000000","0011100100011011","0011000111011000","1111000111000010",
"1100001011110100","1101101000110011","0001111000111000","0011111111111101",
"0001100011000101","1101011011010001","1100001100010010","1111011100111111",
"0011010100100011","0011011011100000","1111101011000001","1100010011101011",
"1101001100101101","0001010100111100","0011111100000110","0010000011001010",
"1101110111001011","1100000100001001","1110111000111101","0010111100101010",
"0011101111101000","0000001111000001","1100100011100010","1100110100100110",
"0000110000111110","0011111000001111","0010100011001111","1110010111000111",
"1100000000000000","1110010100111001","0010100000110001","0011111011110001",
"0000110011000010","1100110111011010","1100100000011110","0000001100111111",
"0011101100011000","0010111111010110","1110111011000011","1100000111110111",
"1101110100110101","0010000000110110","0011111111111010","0001010111000100",
"1101001111010011","1100010000010101","1111101000111111","0011011000100000",
"0011010111011101","1111011111000001","1100001111101110","1101011000101111",
"0001100000111011","0011111100000011","0001111011001000","1101101011001101",
"1100001000001100","1111000100111110","0011000100101000","0011100111100101",
"0000000011000000","1100011111100101","1100111100101000","0000111100111110",
"0011111000001100","0010011011001101","1110001011001000","1100000100000011",
"1110100000111011","0010101000101111","0011110111101110","0000100111000001",
"1100101111011101","1100101000100000","0000011000111111","0011110000010101",
"0010110111010011","1110101111000100","1100000111111010","1110000000110110",
"0010001100110101","0011111111110111","0001001011000011","1101000111010110",
"1100010100011000","1111110100111111","0011100000011110","0011001111011010",
"1111010011000010","1100001011110001","1101100000110001","0001101100111001",
"0100000000000000","1110101111000100","1100111100101000","0011011000100000",
"0000110011000010","1100000100001001","0001111000111000","0010101011010001",
"1100010111101000","1111110100111111","0011110111101110","1101101011001101",
"1101110100110101","0011111000001111","1111101011000001","1100011100011011",
"0010110100101101","0001101111000111","1100000111111010","0000111100111110",
"0011010111011101","1100110111011010","1110111000111101","0011111111111101",
"1110100011000101","1101000100101010","0011100000011110","0000100111000001",
"1100001000001100","0010000000110110","0010100011001111","1100010011101011",
"0000000001000000","0011110011101011","1101100011001111","1110000000110110",
"0011111000001100","1111011111000001","1100100000011110","0010111100101010",
"0001100011000101","1100000111111101","0001001000111101","0011001111011010",
"1100101111011101","1111000100111110","0011111111111010","1110010111000111",
"1101001100101101","0011100100011011","0000011011000001","1100001000001111",
"0010001100110101","0010011011001101","1100001111101110","0000001100111111",
"0011101111101000","1101011011010001","1110001000111000","0011111100001001",
"1111010011000010","1100101000100000","0011000100101000","0001010111000100",
"1100000000000000","0001010100111100","0011000111011000","1100101011100000",
"1111010000111110","0011111111110111","1110001011001000","1101011000101111",
"0011101100011000","0000001111000001","1100001100010010","0010011000110011",
"0010001111001011","1100001011110001","0000011000111111","0011100111100101",
"1101001111010011","1110010100111001","0011111100000110","1111000111000010",
"1100101100100011","0011001100100110","0001001011000011","1100000100000011",
"0001100000111011","0010111111010110","1100100011100010","1111011100111111",
"0011111011110100","1110000011001010","1101100000110001","0011110000010101",
"0000000011000000","1100010000010101","0010100000110001","0010000011001010",
"1100001011110100","0000100100111111","0011100011100010","1101000111010110",
"1110100000111011","0011111100000011","1110111011000011","1100110100100110",
"0011010100100011","0000111111000010","1100000100000110","0001101100111001",
"0010110111010011","1100011111100101","1111101000111111","0011111011110001",
"1101110111001011","1101101000110011","0011110100010010","1111110111000001",
"1100010100011000","0010101000101111","0001111011001000","1100000111110111",
"0000110000111110","0011011011100000","1100111111011000","1110101100111100",
"0100000000000000","1100011111100101","0010100000110001","1111000111000010",
"1111010000111110","0010011011001101","1100100000011110","0011111111111101",
"1100010111101000","0010101000101111","1110111011000011","1111011100111111",
"0010001111001011","1100101000100000","0011111111111010","1100010011101011",
"0010110100101101","1110101111000100","1111101000111111","0010000011001010",
"1100101100100011","0011111111110111","1100001111101110","0010111100101010",
"1110100011000101","1111110100111111","0001111011001000","1100110100100110",
"0011111011110100","1100001011110001","0011000100101000","1110010111000111",
"0000000001000000","0001101111000111","1100111100101000","0011111011110001",
"1100001011110100","0011001100100110","1110001011001000","0000001100111111",
"0001100011000101","1101000100101010","0011110111101110","1100000111110111",
"0011010100100011","1110000011001010","0000011000111111","0001010111000100",
"1101001100101101","0011110011101011","1100000111111010","0011011000100000",
"1101110111001011","0000100100111111","0001001011000011","1101011000101111",
"0011101111101000","1100000111111101","0011100000011110","1101101011001101",
"0000110000111110","0000111111000010","1101100000110001","0011100111100101",
"1100000000000000","0011100100011011","1101100011001111","0000111100111110",
"0000110011000010","1101101000110011","0011100011100010","1100000100000011",
"0011101100011000","1101011011010001","0001001000111101","0000100111000001",
"1101110100110101","0011011011100000","1100000100000110","0011110000010101",
"1101001111010011","0001010100111100","0000011011000001","1110000000110110",
"0011010111011101","1100000100001001","0011110100010010","1101000111010110",
"0001100000111011","0000001111000001","1110001000111000","0011001111011010",
"1100001000001100","0011111000001111","1100111111011000","0001101100111001",
"0000000011000000","1110010100111001","0011000111011000","1100001000001111",
"0011111000001100","1100110111011010","0001111000111000","1111110111000001",
"1110100000111011","0010111111010110","1100001100010010","0011111100001001",
"1100101111011101","0010000000110110","1111101011000001","1110101100111100",
"0010110111010011","1100010000010101","0011111100000110","1100101011100000",
"0010001100110101","1111011111000001","1110111000111101","0010101011010001",
"1100010100011000","0011111100000011","1100100011100010","0010011000110011",
"1111010011000010","1111000100111110","0010100011001111","1100011100011011"
),
("0100000000000000","0011101111101000","0010110111010011","0001100011000101",
"0000000011000000","1110100011000101","1101001111010011","1100010111101000",
"1100000000000000","1100010100011000","1101001100101101","1110100000111011",
"0000000001000000","0001100000111011","0010110100101101","0011101100011000",
"0100000000000000","0011101111101000","0010110111010011","0001100011000101",
"0000000011000000","1110100011000101","1101001111010011","1100010111101000",
"1100000000000000","1100010100011000","1101001100101101","1110100000111011",
"0000000001000000","0001100000111011","0010110100101101","0011101100011000",
"0100000000000000","0011101111101000","0010110111010011","0001100011000101",
"0000000011000000","1110100011000101","1101001111010011","1100010111101000",
"1100000000000000","1100010100011000","1101001100101101","1110100000111011",
"0000000001000000","0001100000111011","0010110100101101","0011101100011000",
"0100000000000000","0011101111101000","0010110111010011","0001100011000101",
"0000000011000000","1110100011000101","1101001111010011","1100010111101000",
"1100000000000000","1100010100011000","1101001100101101","1110100000111011",
"0000000001000000","0001100000111011","0010110100101101","0011101100011000",
"0100000000000000","0011101111101000","0010110111010011","0001100011000101",
"0000000011000000","1110100011000101","1101001111010011","1100010111101000",
"1100000000000000","1100010100011000","1101001100101101","1110100000111011",
"0000000001000000","0001100000111011","0010110100101101","0011101100011000",
"0100000000000000","0011101111101000","0010110111010011","0001100011000101",
"0000000011000000","1110100011000101","1101001111010011","1100010111101000",
"1100000000000000","1100010100011000","1101001100101101","1110100000111011",
"0000000001000000","0001100000111011","0010110100101101","0011101100011000",
"0100000000000000","0011101111101000","0010110111010011","0001100011000101",
"0000000011000000","1110100011000101","1101001111010011","1100010111101000",
"1100000000000000","1100010100011000","1101001100101101","1110100000111011",
"0000000001000000","0001100000111011","0010110100101101","0011101100011000",
"0100000000000000","0011101111101000","0010110111010011","0001100011000101",
"0000000011000000","1110100011000101","1101001111010011","1100010111101000",
"1100000000000000","1100010100011000","1101001100101101","1110100000111011",
"0000000001000000","0001100000111011","0010110100101101","0011101100011000",
"0100000000000000","0001100011000101","1101001111010011","1100010100011000",
"0000000001000000","0011101100011000","0010110111010011","1110100011000101",
"1100000000000000","1110100000111011","0010110100101101","0011101111101000",
"0000000011000000","1100010111101000","1101001100101101","0001100000111011",
"0100000000000000","0001100011000101","1101001111010011","1100010100011000",
"0000000001000000","0011101100011000","0010110111010011","1110100011000101",
"1100000000000000","1110100000111011","0010110100101101","0011101111101000",
"0000000011000000","1100010111101000","1101001100101101","0001100000111011",
"0100000000000000","0001100011000101","1101001111010011","1100010100011000",
"0000000001000000","0011101100011000","0010110111010011","1110100011000101",
"1100000000000000","1110100000111011","0010110100101101","0011101111101000",
"0000000011000000","1100010111101000","1101001100101101","0001100000111011",
"0100000000000000","0001100011000101","1101001111010011","1100010100011000",
"0000000001000000","0011101100011000","0010110111010011","1110100011000101",
"1100000000000000","1110100000111011","0010110100101101","0011101111101000",
"0000000011000000","1100010111101000","1101001100101101","0001100000111011",
"0100000000000000","0001100011000101","1101001111010011","1100010100011000",
"0000000001000000","0011101100011000","0010110111010011","1110100011000101",
"1100000000000000","1110100000111011","0010110100101101","0011101111101000",
"0000000011000000","1100010111101000","1101001100101101","0001100000111011",
"0100000000000000","0001100011000101","1101001111010011","1100010100011000",
"0000000001000000","0011101100011000","0010110111010011","1110100011000101",
"1100000000000000","1110100000111011","0010110100101101","0011101111101000",
"0000000011000000","1100010111101000","1101001100101101","0001100000111011",
"0100000000000000","0001100011000101","1101001111010011","1100010100011000",
"0000000001000000","0011101100011000","0010110111010011","1110100011000101",
"1100000000000000","1110100000111011","0010110100101101","0011101111101000",
"0000000011000000","1100010111101000","1101001100101101","0001100000111011",
"0100000000000000","0001100011000101","1101001111010011","1100010100011000",
"0000000001000000","0011101100011000","0010110111010011","1110100011000101",
"1100000000000000","1110100000111011","0010110100101101","0011101111101000",
"0000000011000000","1100010111101000","1101001100101101","0001100000111011",
"0100000000000000","1110100011000101","1101001100101101","0011101100011000",
"0000000011000000","1100010100011000","0010110100101101","0001100011000101",
"1100000000000000","0001100000111011","0010110111010011","1100010111101000",
"0000000001000000","0011101111101000","1101001111010011","1110100000111011",
"0100000000000000","1110100011000101","1101001100101101","0011101100011000",
"0000000011000000","1100010100011000","0010110100101101","0001100011000101",
"1100000000000000","0001100000111011","0010110111010011","1100010111101000",
"0000000001000000","0011101111101000","1101001111010011","1110100000111011",
"0100000000000000","1110100011000101","1101001100101101","0011101100011000",
"0000000011000000","1100010100011000","0010110100101101","0001100011000101",
"1100000000000000","0001100000111011","0010110111010011","1100010111101000",
"0000000001000000","0011101111101000","1101001111010011","1110100000111011",
"0100000000000000","1110100011000101","1101001100101101","0011101100011000",
"0000000011000000","1100010100011000","0010110100101101","0001100011000101",
"1100000000000000","0001100000111011","0010110111010011","1100010111101000",
"0000000001000000","0011101111101000","1101001111010011","1110100000111011",
"0100000000000000","1110100011000101","1101001100101101","0011101100011000",
"0000000011000000","1100010100011000","0010110100101101","0001100011000101",
"1100000000000000","0001100000111011","0010110111010011","1100010111101000",
"0000000001000000","0011101111101000","1101001111010011","1110100000111011",
"0100000000000000","1110100011000101","1101001100101101","0011101100011000",
"0000000011000000","1100010100011000","0010110100101101","0001100011000101",
"1100000000000000","0001100000111011","0010110111010011","1100010111101000",
"0000000001000000","0011101111101000","1101001111010011","1110100000111011",
"0100000000000000","1110100011000101","1101001100101101","0011101100011000",
"0000000011000000","1100010100011000","0010110100101101","0001100011000101",
"1100000000000000","0001100000111011","0010110111010011","1100010111101000",
"0000000001000000","0011101111101000","1101001111010011","1110100000111011",
"0100000000000000","1110100011000101","1101001100101101","0011101100011000",
"0000000011000000","1100010100011000","0010110100101101","0001100011000101",
"1100000000000000","0001100000111011","0010110111010011","1100010111101000",
"0000000001000000","0011101111101000","1101001111010011","1110100000111011",
"0100000000000000","1100010111101000","0010110100101101","1110100011000101",
"0000000001000000","0001100011000101","1101001100101101","0011101111101000",
"1100000000000000","0011101100011000","1101001111010011","0001100000111011",
"0000000011000000","1110100000111011","0010110111010011","1100010100011000",
"0100000000000000","1100010111101000","0010110100101101","1110100011000101",
"0000000001000000","0001100011000101","1101001100101101","0011101111101000",
"1100000000000000","0011101100011000","1101001111010011","0001100000111011",
"0000000011000000","1110100000111011","0010110111010011","1100010100011000",
"0100000000000000","1100010111101000","0010110100101101","1110100011000101",
"0000000001000000","0001100011000101","1101001100101101","0011101111101000",
"1100000000000000","0011101100011000","1101001111010011","0001100000111011",
"0000000011000000","1110100000111011","0010110111010011","1100010100011000",
"0100000000000000","1100010111101000","0010110100101101","1110100011000101",
"0000000001000000","0001100011000101","1101001100101101","0011101111101000",
"1100000000000000","0011101100011000","1101001111010011","0001100000111011",
"0000000011000000","1110100000111011","0010110111010011","1100010100011000",
"0100000000000000","1100010111101000","0010110100101101","1110100011000101",
"0000000001000000","0001100011000101","1101001100101101","0011101111101000",
"1100000000000000","0011101100011000","1101001111010011","0001100000111011",
"0000000011000000","1110100000111011","0010110111010011","1100010100011000",
"0100000000000000","1100010111101000","0010110100101101","1110100011000101",
"0000000001000000","0001100011000101","1101001100101101","0011101111101000",
"1100000000000000","0011101100011000","1101001111010011","0001100000111011",
"0000000011000000","1110100000111011","0010110111010011","1100010100011000",
"0100000000000000","1100010111101000","0010110100101101","1110100011000101",
"0000000001000000","0001100011000101","1101001100101101","0011101111101000",
"1100000000000000","0011101100011000","1101001111010011","0001100000111011",
"0000000011000000","1110100000111011","0010110111010011","1100010100011000",
"0100000000000000","1100010111101000","0010110100101101","1110100011000101",
"0000000001000000","0001100011000101","1101001100101101","0011101111101000",
"1100000000000000","0011101100011000","1101001111010011","0001100000111011",
"0000000011000000","1110100000111011","0010110111010011","1100010100011000"
),
("0100000000000000","0011100111100101","0010100011001111","0000111111000010",
"1111010011000010","1101101011001101","1100100011100010","1100000111111101",
"1100010100011000","1101011000101111","1110111000111101","0000100100111111",
"0010001100110101","0011011000100000","0011111100000110","0011110011101011",
"0010110111010011","0001010111000100","1111101011000001","1110000011001010",
"1100101111011101","1100000111110111","1100001100010010","1101000100101010",
"1110100000111011","0000001100111111","0001111000111000","0011001100100110",
"0011111000001100","0011111011110001","0011000111011000","0001101111000111",
"0000000011000000","1110010111000111","1100111111011000","1100001011110001",
"1100001000001100","1100110100100110","1110001000111000","1111110100111111",
"0001100000111011","0010111100101010","0011110100010010","0011111111110111",
"0011010111011101","0010000011001010","0000011011000001","1110101111000100",
"1101001111010011","1100010011101011","1100000100000110","1100101000100000",
"1101110100110101","1111011100111111","0001001000111101","0010101000101111",
"0011101100011000","0011111111111101","0011100011100010","0010011011001101",
"0000110011000010","1111000111000010","1101100011001111","1100011111100101",
"1100000000000000","1100011100011011","1101100000110001","1111000100111110",
"0000110000111110","0010011000110011","0011100000011110","0011111100000011",
"0011101111101000","0010101011010001","0001001011000011","1111011111000001",
"1101110111001011","1100101011100000","1100000111111010","1100010000010101",
"1101001100101101","1110101100111100","0000011000111111","0010000000110110",
"0011010100100011","0011111100001001","0011110111101110","0010111111010110",
"0001100011000101","1111110111000001","1110001011001000","1100110111011010",
"1100001011110100","1100001000001111","1100111100101000","1110010100111001",
"0000000001000000","0001101100111001","0011000100101000","0011111000001111",
"0011111011110100","0011001111011010","0001111011001000","0000001111000001",
"1110100011000101","1101000111010110","1100001111101110","1100000100001001",
"1100101100100011","1110000000110110","1111101000111111","0001010100111100",
"0010110100101101","0011110000010101","0011111111111010","0011011011100000",
"0010001111001011","0000100111000001","1110111011000011","1101011011010001",
"1100010111101000","1100000100000011","1100100000011110","1101101000110011",
"1111010000111110","0000111100111110","0010100000110001","0011100100011011",
"0100000000000000","0001010111000100","1100111111011000","1100101000100000",
"0000110000111110","0011111100001001","0001111011001000","1101011011010001",
"1100010100011000","0000001100111111","0011110100010010","0010011011001101",
"1101110111001011","1100001000001111","1111101000111111","0011100100011011",
"0010110111010011","1110010111000111","1100000100000110","1111000100111110",
"0011010100100011","0011001111011010","1110111011000011","1100000111111101",
"1110100000111011","0010111100101010","0011100011100010","1111011111000001",
"1100001011110100","1110000000110110","0010100000110001","0011110011101011",
"0000000011000000","1100010011101011","1101100000110001","0010000000110110",
"0011111011110100","0000100111000001","1100100011100010","1101000100101010",
"0001100000111011","0011111111111101","0001001011000011","1100110111011010",
"1100101100100011","0000111100111110","0011111100000110","0001101111000111",
"1101001111010011","1100011100011011","0000011000111111","0011111000001111",
"0010001111001011","1101101011001101","1100001100010010","1111110100111111",
"0011101100011000","0010101011010001","1110001011001000","1100000100001001",
"1111010000111110","0011011000100000","0011000111011000","1110101111000100",
"1100000000000000","1110101100111100","0011000100101000","0011011011100000",
"1111010011000010","1100000111110111","1110001000111000","0010101000101111",
"0011101111101000","1111110111000001","1100001111101110","1101101000110011",
"0010001100110101","0011111011110001","0000011011000001","1100011111100101",
"1101001100101101","0001101100111001","0011111111111010","0000111111000010",
"1100101111011101","1100110100100110","0001001000111101","0011111100000011",
"0001100011000101","1101000111010110","1100100000011110","0000100100111111",
"0011111000001100","0010000011001010","1101100011001111","1100010000010101",
"0000000001000000","0011110000010101","0010100011001111","1110000011001010",
"1100001000001100","1111011100111111","0011100000011110","0010111111010110",
"1110100011000101","1100000100000011","1110111000111101","0011001100100110",
"0011010111011101","1111000111000010","1100000111111010","1110010100111001",
"0010110100101101","0011100111100101","1111101011000001","1100001011110001",
"1101110100110101","0010011000110011","0011110111101110","0000001111000001",
"1100010111101000","1101011000101111","0001111000111000","0011111111110111",
"0000110011000010","1100101011100000","1100111100101000","0001010100111100",
"0100000000000000","1110010111000111","1101100000110001","0011111000001111",
"1111010011000010","1100110100100110","0011100000011110","0000001111000001",
"1100010100011000","0010111100101010","0001001011000011","1100000100001001",
"0010001100110101","0010000011001010","1100000111111010","0001010100111100",
"0010110111010011","1100010011101011","0000011000111111","0011011011100000",
"1100101111011101","1111011100111111","0011110111101110","1101011011010001",
"1110100000111011","0011111111111101","1110001011001000","1101101000110011",
"0011111000001100","1111000111000010","1100111100101000","0011100100011011",
"0000000011000000","1100011100011011","0011000100101000","0000111111000010",
"1100001000001100","0010011000110011","0001111011001000","1100000111111101",
"0001100000111011","0010101011010001","1100001111101110","0000100100111111",
"0011010111011101","1100101011100000","1111101000111111","0011110011101011",
"1101001111010011","1110101100111100","0011111111111010","1110000011001010",
"1101110100110101","0011111100001001","1110111011000011","1101000100101010",
"0011101100011000","1111110111000001","1100100000011110","0011001100100110",
"0000110011000010","1100001000001111","0010100000110001","0001101111000111",
"1100000000000000","0001101100111001","0010100011001111","1100001011110001",
"0000110000111110","0011001111011010","1100100011100010","1111110100111111",
"0011101111101000","1101000111010110","1110111000111101","0011111111110111",
"1101110111001011","1110000000110110","0011111100000110","1110101111000100",
"1101001100101101","0011110000010101","1111101011000001","1100101000100000",
"0011010100100011","0000100111000001","1100001100010010","0010101000101111",
"0001100011000101","1100000100000011","0001111000111000","0010011011001101",
"1100001011110100","0000111100111110","0011000111011000","1100011111100101",
"0000000001000000","0011100111100101","1100111111011000","1111000100111110",
"0011111011110100","1101101011001101","1110001000111000","0011111100000011",
"1110100011000101","1101011000101111","0011110100010010","1111011111000001",
"1100101100100011","0011011000100000","0000011011000001","1100010000010101",
"0010110100101101","0001010111000100","1100000100000110","0010000000110110",
"0010001111001011","1100000111110111","0001001000111101","0010111111010110",
"1100010111101000","0000001100111111","0011100011100010","1100110111011010",
"1111010000111110","0011111011110001","1101100011001111","1110010100111001",
"0100000000000000","1100010011101011","0011000100101000","1110000011001010",
"0000110000111110","0000100111000001","1110001000111000","0010111111010110",
"1100010100011000","0011111111111101","1100001111101110","0011001100100110",
"1101110111001011","0000111100111110","0000011011000001","1110010100111001",
"0010110111010011","1100011100011011","0011111111111010","1100001011110001",
"0011010100100011","1101101011001101","0001001000111101","0000001111000001",
"1110100000111011","0010101011010001","1100100000011110","0011111111110111",
"1100001011110100","0011011000100000","1101100011001111","0001010100111100",
"0000000011000000","1110101100111100","0010100011001111","1100101000100000",
"0011111011110100","1100000111110111","0011100000011110","1101011011010001",
"0001100000111011","1111110111000001","1110111000111101","0010011011001101",
"1100101100100011","0011111011110001","1100000111111010","0011100100011011",
"1101001111010011","0001101100111001","1111101011000001","1111000100111110",
"0010001111001011","1100110100100110","0011110111101110","1100000111111101",
"0011101100011000","1101000111010110","0001111000111000","1111011111000001",
"1111010000111110","0010000011001010","1100111100101000","0011110011101011",
"1100000000000000","0011110000010101","1100111111011000","0010000000110110",
"1111010011000010","1111011100111111","0001111011001000","1101000100101010",
"0011101111101000","1100000100000011","0011110100010010","1100110111011010",
"0010001100110101","1111000111000010","1111101000111111","0001101111000111",
"1101001100101101","0011100111100101","1100000100000110","0011111000001111",
"1100101111011101","0010011000110011","1110111011000011","1111110100111111",
"0001100011000101","1101011000101111","0011100011100010","1100000100001001",
"0011111000001100","1100101011100000","0010100000110001","1110101111000100",
"0000000001000000","0001010111000100","1101100000110001","0011011011100000",
"1100001000001100","0011111100001001","1100100011100010","0010101000101111",
"1110100011000101","0000001100111111","0001001011000011","1101101000110011",
"0011010111011101","1100001000001111","0011111100000110","1100011111100101",
"0010110100101101","1110010111000111","0000011000111111","0000111111000010",
"1101110100110101","0011001111011010","1100001100010010","0011111100000011",
"1100010111101000","0010111100101010","1110001011001000","0000100100111111",
"0000110011000010","1110000000110110","0011000111011000","1100010000010101"
),
("0100000000000000","0011100011100010","0010001111001011","0000011011000001",
"1110100011000101","1100111111011000","1100001011110100","1100001100010010",
"1101001100101101","1110111000111101","0000110000111110","0010100000110001",
"0011101100011000","0011111111111010","0011010111011101","0001111011001000",
"0000000011000000","1110001011001000","1100101111011101","1100000111111010",
"1100010100011000","1101100000110001","1111010000111110","0001001000111101",
"0010110100101101","0011110100010010","0011111011110100","0011000111011000",
"0001100011000101","1111101011000001","1101110111001011","1100100011100010",
"1100000000000000","1100100000011110","1101110100110101","1111101000111111",
"0001100000111011","0011000100101000","0011111000001100","0011110111101110",
"0010110111010011","0001001011000011","1111010011000010","1101100011001111",
"1100010111101000","1100000100000110","1100101100100011","1110001000111000",
"0000000001000000","0001111000111000","0011010100100011","0011111100000110",
"0011101111101000","0010100011001111","0000110011000010","1110111011000011",
"1101001111010011","1100001111101110","1100001000001100","1100111100101000",
"1110100000111011","0000011000111111","0010001100110101","0011100000011110",
"0100000000000000","0011100011100010","0010001111001011","0000011011000001",
"1110100011000101","1100111111011000","1100001011110100","1100001100010010",
"1101001100101101","1110111000111101","0000110000111110","0010100000110001",
"0011101100011000","0011111111111010","0011010111011101","0001111011001000",
"0000000011000000","1110001011001000","1100101111011101","1100000111111010",
"1100010100011000","1101100000110001","1111010000111110","0001001000111101",
"0010110100101101","0011110100010010","0011111011110100","0011000111011000",
"0001100011000101","1111101011000001","1101110111001011","1100100011100010",
"1100000000000000","1100100000011110","1101110100110101","1111101000111111",
"0001100000111011","0011000100101000","0011111000001100","0011110111101110",
"0010110111010011","0001001011000011","1111010011000010","1101100011001111",
"1100010111101000","1100000100000110","1100101100100011","1110001000111000",
"0000000001000000","0001111000111000","0011010100100011","0011111100000110",
"0011101111101000","0010100011001111","0000110011000010","1110111011000011",
"1101001111010011","1100001111101110","1100001000001100","1100111100101000",
"1110100000111011","0000011000111111","0010001100110101","0011100000011110",
"0100000000000000","0001001011000011","1100101111011101","1100111100101000",
"0001100000111011","0011111111111010","0000110011000010","1100100011100010",
"1101001100101101","0001111000111000","0011111011110100","0000011011000001",
"1100010111101000","1101100000110001","0010001100110101","0011110111101110",
"0000000011000000","1100001111101110","1101110100110101","0010100000110001",
"0011101111101000","1111101011000001","1100001011110100","1110001000111000",
"0010110100101101","0011100011100010","1111010011000010","1100000111111010",
"1110100000111011","0011000100101000","0011010111011101","1110111011000011",
"1100000000000000","1110111000111101","0011010100100011","0011000111011000",
"1110100011000101","1100000100000110","1111010000111110","0011100000011110",
"0010110111010011","1110001011001000","1100001000001100","1111101000111111",
"0011101100011000","0010100011001111","1101110111001011","1100001100010010",
"0000000001000000","0011110100010010","0010001111001011","1101100011001111",
"1100010100011000","0000011000111111","0011111000001100","0001111011001000",
"1101001111010011","1100100000011110","0000110000111110","0011111100000110",
"0001100011000101","1100111111011000","1100101100100011","0001001000111101",
"0100000000000000","0001001011000011","1100101111011101","1100111100101000",
"0001100000111011","0011111111111010","0000110011000010","1100100011100010",
"1101001100101101","0001111000111000","0011111011110100","0000011011000001",
"1100010111101000","1101100000110001","0010001100110101","0011110111101110",
"0000000011000000","1100001111101110","1101110100110101","0010100000110001",
"0011101111101000","1111101011000001","1100001011110100","1110001000111000",
"0010110100101101","0011100011100010","1111010011000010","1100000111111010",
"1110100000111011","0011000100101000","0011010111011101","1110111011000011",
"1100000000000000","1110111000111101","0011010100100011","0011000111011000",
"1110100011000101","1100000100000110","1111010000111110","0011100000011110",
"0010110111010011","1110001011001000","1100001000001100","1111101000111111",
"0011101100011000","0010100011001111","1101110111001011","1100001100010010",
"0000000001000000","0011110100010010","0010001111001011","1101100011001111",
"1100010100011000","0000011000111111","0011111000001100","0001111011001000",
"1101001111010011","1100100000011110","0000110000111110","0011111100000110",
"0001100011000101","1100111111011000","1100101100100011","0001001000111101",
"0100000000000000","1110001011001000","1101110100110101","0011111100000110",
"1110100011000101","1101100000110001","0011111000001100","1110111011000011",
"1101001100101101","0011110100010010","1111010011000010","1100111100101000",
"0011101100011000","1111101011000001","1100101100100011","0011100000011110",
"0000000011000000","1100100000011110","0011010100100011","0000011011000001",
"1100010100011000","0011000100101000","0000110011000010","1100001100010010",
"0010110100101101","0001001011000011","1100001000001100","0010100000110001",
"0001100011000101","1100000100000110","0010001100110101","0001111011001000",
"1100000000000000","0001111000111000","0010001111001011","1100000111111010",
"0001100000111011","0010100011001111","1100001011110100","0001001000111101",
"0010110111010011","1100001111101110","0000110000111110","0011000111011000",
"1100010111101000","0000011000111111","0011010111011101","1100100011100010",
"0000000001000000","0011100011100010","1100101111011101","1111101000111111",
"0011101111101000","1100111111011000","1111010000111110","0011110111101110",
"1101001111010011","1110111000111101","0011111011110100","1101100011001111",
"1110100000111011","0011111111111010","1101110111001011","1110001000111000",
"0100000000000000","1110001011001000","1101110100110101","0011111100000110",
"1110100011000101","1101100000110001","0011111000001100","1110111011000011",
"1101001100101101","0011110100010010","1111010011000010","1100111100101000",
"0011101100011000","1111101011000001","1100101100100011","0011100000011110",
"0000000011000000","1100100000011110","0011010100100011","0000011011000001",
"1100010100011000","0011000100101000","0000110011000010","1100001100010010",
"0010110100101101","0001001011000011","1100001000001100","0010100000110001",
"0001100011000101","1100000100000110","0010001100110101","0001111011001000",
"1100000000000000","0001111000111000","0010001111001011","1100000111111010",
"0001100000111011","0010100011001111","1100001011110100","0001001000111101",
"0010110111010011","1100001111101110","0000110000111110","0011000111011000",
"1100010111101000","0000011000111111","0011010111011101","1100100011100010",
"0000000001000000","0011100011100010","1100101111011101","1111101000111111",
"0011101111101000","1100111111011000","1111010000111110","0011110111101110",
"1101001111010011","1110111000111101","0011111011110100","1101100011001111",
"1110100000111011","0011111111111010","1101110111001011","1110001000111000",
"0100000000000000","1100001111101110","0011010100100011","1101100011001111",
"0001100000111011","1111101011000001","1111010000111110","0001111011001000",
"1101001100101101","0011100011100010","1100001000001100","0011111100000110",
"1100010111101000","0011000100101000","1101110111001011","0001001000111101",
"0000000011000000","1110111000111101","0010001111001011","1100111100101000",
"0011101111101000","1100000100000110","0011111000001100","1100100011100010",
"0010110100101101","1110001011001000","0000110000111110","0000011011000001",
"1110100000111011","0010100011001111","1100101100100011","0011110111101110",
"1100000000000000","0011110100010010","1100101111011101","0010100000110001",
"1110100011000101","0000011000111111","0000110011000010","1110001000111000",
"0010110111010011","1100100000011110","0011111011110100","1100000111111010",
"0011101100011000","1100111111011000","0010001100110101","1110111011000011",
"0000000001000000","0001001011000011","1101110100110101","0011000111011000",
"1100010100011000","0011111111111010","1100001011110100","0011100000011110",
"1101001111010011","0001111000111000","1111010011000010","1111101000111111",
"0001100011000101","1101100000110001","0011010111011101","1100001100010010",
"0100000000000000","1100001111101110","0011010100100011","1101100011001111",
"0001100000111011","1111101011000001","1111010000111110","0001111011001000",
"1101001100101101","0011100011100010","1100001000001100","0011111100000110",
"1100010111101000","0011000100101000","1101110111001011","0001001000111101",
"0000000011000000","1110111000111101","0010001111001011","1100111100101000",
"0011101111101000","1100000100000110","0011111000001100","1100100011100010",
"0010110100101101","1110001011001000","0000110000111110","0000011011000001",
"1110100000111011","0010100011001111","1100101100100011","0011110111101110",
"1100000000000000","0011110100010010","1100101111011101","0010100000110001",
"1110100011000101","0000011000111111","0000110011000010","1110001000111000",
"0010110111010011","1100100000011110","0011111011110100","1100000111111010",
"0011101100011000","1100111111011000","0010001100110101","1110111011000011",
"0000000001000000","0001001011000011","1101110100110101","0011000111011000",
"1100010100011000","0011111111111010","1100001011110100","0011100000011110",
"1101001111010011","0001111000111000","1111010011000010","1111101000111111",
"0001100011000101","1101100000110001","0011010111011101","1100001100010010"
),
("0100000000000000","0011011011100000","0001111011001000","1111110111000001",
"1101110111001011","1100011111100101","1100000100000110","1100110100100110",
"1110100000111011","0000100100111111","0010100000110001","0011110000010101",
"0011111011110100","0010111111010110","0001001011000011","1111000111000010",
"1101001111010011","1100001011110001","1100001100010010","1101011000101111",
"1111010000111110","0001010100111100","0011000100101000","0011111100001001",
"0011101111101000","0010011011001101","0000011011000001","1110010111000111",
"1100101111011101","1100000111111101","1100100000011110","1110000000110110",
"0000000001000000","0010000000110110","0011100000011110","0011111111111101",
"0011010111011101","0001101111000111","1111101011000001","1101101011001101",
"1100010111101000","1100000100001001","1100111100101000","1110101100111100",
"0000110000111110","0010101000101111","0011110100010010","0011111011110001",
"0010110111010011","0000111111000010","1110111011000011","1101000111010110",
"1100001011110100","1100010000010101","1101100000110001","1111011100111111",
"0001100000111011","0011001100100110","0011111100000110","0011100111100101",
"0010001111001011","0000001111000001","1110001011001000","1100101011100000",
"1100000000000000","1100101000100000","1110001000111000","0000001100111111",
"0010001100110101","0011100100011011","0011111111111010","0011001111011010",
"0001100011000101","1111011111000001","1101100011001111","1100010011101011",
"1100001000001100","1101000100101010","1110111000111101","0000111100111110",
"0010110100101101","0011111000001111","0011110111101110","0010101011010001",
"0000110011000010","1110101111000100","1100111111011000","1100000111110111",
"1100010100011000","1101101000110011","1111101000111111","0001101100111001",
"0011010100100011","0011111100000011","0011100011100010","0010000011001010",
"0000000011000000","1110000011001010","1100100011100010","1100000100000011",
"1100101100100011","1110010100111001","0000011000111111","0010011000110011",
"0011101100011000","0011111111110111","0011000111011000","0001010111000100",
"1111010011000010","1101011011010001","1100001111101110","1100001000001111",
"1101001100101101","1111000100111110","0001001000111101","0010111100101010",
"0011111000001100","0011110011101011","0010100011001111","0000100111000001",
"1110100011000101","1100110111011010","1100000111111010","1100011100011011",
"1101110100110101","1111110100111111","0001111000111000","0011011000100000",
"0100000000000000","0000111111000010","1100100011100010","1101011000101111",
"0010001100110101","0011110011101011","1111101011000001","1100000111110111",
"1110100000111011","0011001100100110","0011000111011000","1110010111000111",
"1100001000001100","1111110100111111","0011110100010010","0010000011001010",
"1101001111010011","1100101000100000","0001001000111101","0011111111111101",
"0000110011000010","1100011111100101","1101100000110001","0010011000110011",
"0011101111101000","1111011111000001","1100000111111010","1110101100111100",
"0011010100100011","0010111111010110","1110001011001000","1100001000001111",
"0000000001000000","0011111000001111","0001111011001000","1101000111010110",
"1100101100100011","0001010100111100","0011111111111010","0000100111000001",
"1100010111101000","1101101000110011","0010100000110001","0011100111100101",
"1111010011000010","1100000111111101","1110111000111101","0011011000100000",
"0010110111010011","1110000011001010","1100001100010010","0000001100111111",
"0011111000001100","0001101111000111","1100111111011000","1100110100100110",
"0001100000111011","0011111111110111","0000011011000001","1100010011101011",
"1101110100110101","0010101000101111","0011100011100010","1111000111000010",
"1100000000000000","1111000100111110","0011100000011110","0010101011010001",
"1101110111001011","1100010000010101","0000011000111111","0011111100001001",
"0001100011000101","1100110111011010","1100111100101000","0001101100111001",
"0011111011110100","0000001111000001","1100001111101110","1110000000110110",
"0010110100101101","0011011011100000","1110111011000011","1100000100000011",
"1111010000111110","0011100100011011","0010100011001111","1101101011001101",
"1100010100011000","0000100100111111","0011111100000110","0001010111000100",
"1100101111011101","1101000100101010","0001111000111000","0011111011110001",
"0000000011000000","1100001011110001","1110001000111000","0010111100101010",
"0011010111011101","1110101111000100","1100000100000110","1111011100111111",
"0011101100011000","0010011011001101","1101100011001111","1100011100011011",
"0000110000111110","0011111100000011","0001001011000011","1100101011100000",
"1101001100101101","0010000000110110","0011110111101110","1111110111000001",
"1100001011110100","1110010100111001","0011000100101000","0011001111011010",
"1110100011000101","1100000100001001","1111101000111111","0011110000010101",
"0010001111001011","1101011011010001","1100100000011110","0000111100111110",
"0100000000000000","1110000011001010","1110001000111000","0011111111111101",
"1101110111001011","1110010100111001","0011111111111010","1101101011001101",
"1110100000111011","0011111111110111","1101100011001111","1110101100111100",
"0011111011110100","1101011011010001","1110111000111101","0011111011110001",
"1101001111010011","1111000100111110","0011110111101110","1101000111010110",
"1111010000111110","0011110011101011","1100111111011000","1111011100111111",
"0011101111101000","1100110111011010","1111101000111111","0011100111100101",
"1100101111011101","1111110100111111","0011100011100010","1100101011100000",
"0000000001000000","0011011011100000","1100100011100010","0000001100111111",
"0011010111011101","1100011111100101","0000011000111111","0011001111011010",
"1100010111101000","0000100100111111","0011000111011000","1100010011101011",
"0000110000111110","0010111111010110","1100001111101110","0000111100111110",
"0010110111010011","1100001011110001","0001001000111101","0010101011010001",
"1100001011110100","0001010100111100","0010100011001111","1100000111110111",
"0001100000111011","0010011011001101","1100000111111010","0001101100111001",
"0010001111001011","1100000111111101","0001111000111000","0010000011001010",
"1100000000000000","0010000000110110","0001111011001000","1100000100000011",
"0010001100110101","0001101111000111","1100000100000110","0010011000110011",
"0001100011000101","1100000100001001","0010100000110001","0001010111000100",
"1100001000001100","0010101000101111","0001001011000011","1100001000001111",
"0010110100101101","0000111111000010","1100001100010010","0010111100101010",
"0000110011000010","1100010000010101","0011000100101000","0000100111000001",
"1100010100011000","0011001100100110","0000011011000001","1100011100011011",
"0011010100100011","0000001111000001","1100100000011110","0011011000100000",
"0000000011000000","1100101000100000","0011100000011110","1111110111000001",
"1100101100100011","0011100100011011","1111101011000001","1100110100100110",
"0011101100011000","1111011111000001","1100111100101000","0011110000010101",
"1111010011000010","1101000100101010","0011110100010010","1111000111000010",
"1101001100101101","0011111000001111","1110111011000011","1101011000101111",
"0011111000001100","1110101111000100","1101100000110001","0011111100001001",
"1110100011000101","1101101000110011","0011111100000110","1110010111000111",
"1101110100110101","0011111100000011","1110001011001000","1110000000110110",
"0100000000000000","1100001011110001","0011100000011110","1101000111010110",
"0010001100110101","1110101111000100","0000011000111111","0000100111000001",
"1110100000111011","0010011011001101","1100111100101000","0011100111100101",
"1100001000001100","0011111100000011","1100001111101110","0011011000100000",
"1101001111010011","0010000000110110","1110111011000011","0000001100111111",
"0000110011000010","1110010100111001","0010100011001111","1100110100100110",
"0011101111101000","1100000100001001","0011111100000110","1100010011101011",
"0011010100100011","1101011011010001","0001111000111000","1111000111000010",
"0000000001000000","0000111111000010","1110001000111000","0010101011010001",
"1100101100100011","0011110011101011","1100000100000110","0011111100001001",
"1100010111101000","0011001100100110","1101100011001111","0001101100111001",
"1111010011000010","1111110100111111","0001001011000011","1110000000110110",
"0010110111010011","1100101000100000","0011110111101110","1100000100000011",
"0011111000001100","1100011111100101","0011000100101000","1101101011001101",
"0001100000111011","1111011111000001","1111101000111111","0001010111000100",
"1101110100110101","0010111111010110","1100100000011110","0011111011110001",
"1100000000000000","0011111000001111","1100100011100010","0010111100101010",
"1101110111001011","0001010100111100","1111101011000001","1111011100111111",
"0001100011000101","1101101000110011","0011000111011000","1100011100011011",
"0011111011110100","1100000111111101","0011110100010010","1100101011100000",
"0010110100101101","1110000011001010","0001001000111101","1111110111000001",
"1111010000111110","0001101111000111","1101100000110001","0011001111011010",
"1100010100011000","0011111111110111","1100000111111010","0011110000010101",
"1100101111011101","0010101000101111","1110001011001000","0000111100111110",
"0000000011000000","1111000100111110","0001111011001000","1101011000101111",
"0011010111011101","1100010000010101","0011111111111010","1100000111110111",
"0011101100011000","1100110111011010","0010100000110001","1110010111000111",
"0000110000111110","0000001111000001","1110111000111101","0010000011001010",
"1101001100101101","0011011011100000","1100001100010010","0011111111111101",
"1100001011110100","0011100100011011","1100111111011000","0010011000110011",
"1110100011000101","0000100100111111","0000011011000001","1110101100111100",
"0010001111001011","1101000100101010","0011100011100010","1100001000001111"
),
("0100000000000000","0011010111011101","0001100011000101","1111010011000010",
"1101001111010011","1100001011110100","1100010100011000","1101110100110101",
"0000000001000000","0010001100110101","0011101100011000","0011111011110100",
"0010110111010011","0000110011000010","1110100011000101","1100101111011101",
"1100000000000000","1100101100100011","1110100000111011","0000110000111110",
"0010110100101101","0011111000001100","0011101111101000","0010001111001011",
"0000000011000000","1101110111001011","1100010111101000","1100001000001100",
"1101001100101101","1111010000111110","0001100000111011","0011010100100011",
"0100000000000000","0011010111011101","0001100011000101","1111010011000010",
"1101001111010011","1100001011110100","1100010100011000","1101110100110101",
"0000000001000000","0010001100110101","0011101100011000","0011111011110100",
"0010110111010011","0000110011000010","1110100011000101","1100101111011101",
"1100000000000000","1100101100100011","1110100000111011","0000110000111110",
"0010110100101101","0011111000001100","0011101111101000","0010001111001011",
"0000000011000000","1101110111001011","1100010111101000","1100001000001100",
"1101001100101101","1111010000111110","0001100000111011","0011010100100011",
"0100000000000000","0011010111011101","0001100011000101","1111010011000010",
"1101001111010011","1100001011110100","1100010100011000","1101110100110101",
"0000000001000000","0010001100110101","0011101100011000","0011111011110100",
"0010110111010011","0000110011000010","1110100011000101","1100101111011101",
"1100000000000000","1100101100100011","1110100000111011","0000110000111110",
"0010110100101101","0011111000001100","0011101111101000","0010001111001011",
"0000000011000000","1101110111001011","1100010111101000","1100001000001100",
"1101001100101101","1111010000111110","0001100000111011","0011010100100011",
"0100000000000000","0011010111011101","0001100011000101","1111010011000010",
"1101001111010011","1100001011110100","1100010100011000","1101110100110101",
"0000000001000000","0010001100110101","0011101100011000","0011111011110100",
"0010110111010011","0000110011000010","1110100011000101","1100101111011101",
"1100000000000000","1100101100100011","1110100000111011","0000110000111110",
"0010110100101101","0011111000001100","0011101111101000","0010001111001011",
"0000000011000000","1101110111001011","1100010111101000","1100001000001100",
"1101001100101101","1111010000111110","0001100000111011","0011010100100011",
"0100000000000000","0000110011000010","1100010111101000","1101110100110101",
"0010110100101101","0011010111011101","1110100011000101","1100001000001100",
"0000000001000000","0011111000001100","0001100011000101","1100101111011101",
"1101001100101101","0010001100110101","0011101111101000","1111010011000010",
"1100000000000000","1111010000111110","0011101100011000","0010001111001011",
"1101001111010011","1100101100100011","0001100000111011","0011111011110100",
"0000000011000000","1100001011110100","1110100000111011","0011010100100011",
"0010110111010011","1101110111001011","1100010100011000","0000110000111110",
"0100000000000000","0000110011000010","1100010111101000","1101110100110101",
"0010110100101101","0011010111011101","1110100011000101","1100001000001100",
"0000000001000000","0011111000001100","0001100011000101","1100101111011101",
"1101001100101101","0010001100110101","0011101111101000","1111010011000010",
"1100000000000000","1111010000111110","0011101100011000","0010001111001011",
"1101001111010011","1100101100100011","0001100000111011","0011111011110100",
"0000000011000000","1100001011110100","1110100000111011","0011010100100011",
"0010110111010011","1101110111001011","1100010100011000","0000110000111110",
"0100000000000000","0000110011000010","1100010111101000","1101110100110101",
"0010110100101101","0011010111011101","1110100011000101","1100001000001100",
"0000000001000000","0011111000001100","0001100011000101","1100101111011101",
"1101001100101101","0010001100110101","0011101111101000","1111010011000010",
"1100000000000000","1111010000111110","0011101100011000","0010001111001011",
"1101001111010011","1100101100100011","0001100000111011","0011111011110100",
"0000000011000000","1100001011110100","1110100000111011","0011010100100011",
"0010110111010011","1101110111001011","1100010100011000","0000110000111110",
"0100000000000000","0000110011000010","1100010111101000","1101110100110101",
"0010110100101101","0011010111011101","1110100011000101","1100001000001100",
"0000000001000000","0011111000001100","0001100011000101","1100101111011101",
"1101001100101101","0010001100110101","0011101111101000","1111010011000010",
"1100000000000000","1111010000111110","0011101100011000","0010001111001011",
"1101001111010011","1100101100100011","0001100000111011","0011111011110100",
"0000000011000000","1100001011110100","1110100000111011","0011010100100011",
"0010110111010011","1101110111001011","1100010100011000","0000110000111110",
"0100000000000000","1101110111001011","1110100000111011","0011111011110100",
"1101001111010011","1111010000111110","0011101111101000","1100101111011101",
"0000000001000000","0011010111011101","1100010111101000","0000110000111110",
"0010110111010011","1100001011110100","0001100000111011","0010001111001011",
"1100000000000000","0010001100110101","0001100011000101","1100001000001100",
"0010110100101101","0000110011000010","1100010100011000","0011010100100011",
"0000000011000000","1100101100100011","0011101100011000","1111010011000010",
"1101001100101101","0011111000001100","1110100011000101","1101110100110101",
"0100000000000000","1101110111001011","1110100000111011","0011111011110100",
"1101001111010011","1111010000111110","0011101111101000","1100101111011101",
"0000000001000000","0011010111011101","1100010111101000","0000110000111110",
"0010110111010011","1100001011110100","0001100000111011","0010001111001011",
"1100000000000000","0010001100110101","0001100011000101","1100001000001100",
"0010110100101101","0000110011000010","1100010100011000","0011010100100011",
"0000000011000000","1100101100100011","0011101100011000","1111010011000010",
"1101001100101101","0011111000001100","1110100011000101","1101110100110101",
"0100000000000000","1101110111001011","1110100000111011","0011111011110100",
"1101001111010011","1111010000111110","0011101111101000","1100101111011101",
"0000000001000000","0011010111011101","1100010111101000","0000110000111110",
"0010110111010011","1100001011110100","0001100000111011","0010001111001011",
"1100000000000000","0010001100110101","0001100011000101","1100001000001100",
"0010110100101101","0000110011000010","1100010100011000","0011010100100011",
"0000000011000000","1100101100100011","0011101100011000","1111010011000010",
"1101001100101101","0011111000001100","1110100011000101","1101110100110101",
"0100000000000000","1101110111001011","1110100000111011","0011111011110100",
"1101001111010011","1111010000111110","0011101111101000","1100101111011101",
"0000000001000000","0011010111011101","1100010111101000","0000110000111110",
"0010110111010011","1100001011110100","0001100000111011","0010001111001011",
"1100000000000000","0010001100110101","0001100011000101","1100001000001100",
"0010110100101101","0000110011000010","1100010100011000","0011010100100011",
"0000000011000000","1100101100100011","0011101100011000","1111010011000010",
"1101001100101101","0011111000001100","1110100011000101","1101110100110101",
"0100000000000000","1100001011110100","0011101100011000","1100101111011101",
"0010110100101101","1101110111001011","0001100000111011","1111010011000010",
"0000000001000000","0000110011000010","1110100000111011","0010001111001011",
"1101001100101101","0011010111011101","1100010100011000","0011111011110100",
"1100000000000000","0011111000001100","1100010111101000","0011010100100011",
"1101001111010011","0010001100110101","1110100011000101","0000110000111110",
"0000000011000000","1111010000111110","0001100011000101","1101110100110101",
"0010110111010011","1100101100100011","0011101111101000","1100001000001100",
"0100000000000000","1100001011110100","0011101100011000","1100101111011101",
"0010110100101101","1101110111001011","0001100000111011","1111010011000010",
"0000000001000000","0000110011000010","1110100000111011","0010001111001011",
"1101001100101101","0011010111011101","1100010100011000","0011111011110100",
"1100000000000000","0011111000001100","1100010111101000","0011010100100011",
"1101001111010011","0010001100110101","1110100011000101","0000110000111110",
"0000000011000000","1111010000111110","0001100011000101","1101110100110101",
"0010110111010011","1100101100100011","0011101111101000","1100001000001100",
"0100000000000000","1100001011110100","0011101100011000","1100101111011101",
"0010110100101101","1101110111001011","0001100000111011","1111010011000010",
"0000000001000000","0000110011000010","1110100000111011","0010001111001011",
"1101001100101101","0011010111011101","1100010100011000","0011111011110100",
"1100000000000000","0011111000001100","1100010111101000","0011010100100011",
"1101001111010011","0010001100110101","1110100011000101","0000110000111110",
"0000000011000000","1111010000111110","0001100011000101","1101110100110101",
"0010110111010011","1100101100100011","0011101111101000","1100001000001100",
"0100000000000000","1100001011110100","0011101100011000","1100101111011101",
"0010110100101101","1101110111001011","0001100000111011","1111010011000010",
"0000000001000000","0000110011000010","1110100000111011","0010001111001011",
"1101001100101101","0011010111011101","1100010100011000","0011111011110100",
"1100000000000000","0011111000001100","1100010111101000","0011010100100011",
"1101001111010011","0010001100110101","1110100011000101","0000110000111110",
"0000000011000000","1111010000111110","0001100011000101","1101110100110101",
"0010110111010011","1100101100100011","0011101111101000","1100001000001100"
),
("0100000000000000","0011001111011010","0001001011000011","1110101111000100",
"1100101111011101","1100000100000011","1100111100101000","1111000100111110",
"0001100000111011","0011011000100000","0011111111111010","0010111111010110",
"0000110011000010","1110010111000111","1100100011100010","1100000100001001",
"1101001100101101","1111011100111111","0001111000111000","0011100100011011",
"0011111011110100","0010101011010001","0000011011000001","1110000011001010",
"1100010111101000","1100001000001111","1101100000110001","1111110100111111",
"0010001100110101","0011110000010101","0011110111101110","0010011011001101",
"0000000011000000","1101101011001101","1100001111101110","1100010000010101",
"1101110100110101","0000001100111111","0010100000110001","0011111000001111",
"0011101111101000","0010000011001010","1111101011000001","1101011011010001",
"1100001011110100","1100011100011011","1110001000111000","0000100100111111",
"0010110100101101","0011111100001001","0011100011100010","0001101111000111",
"1111010011000010","1101000111010110","1100000111111010","1100101000100000",
"1110100000111011","0000111100111110","0011000100101000","0011111100000011",
"0011010111011101","0001010111000100","1110111011000011","1100110111011010",
"1100000000000000","1100110100100110","1110111000111101","0001010100111100",
"0011010100100011","0011111111111101","0011000111011000","0000111111000010",
"1110100011000101","1100101011100000","1100000100000110","1101000100101010",
"1111010000111110","0001101100111001","0011100000011110","0011111111110111",
"0010110111010011","0000100111000001","1110001011001000","1100011111100101",
"1100001000001100","1101011000101111","1111101000111111","0010000000110110",
"0011101100011000","0011111011110001","0010100011001111","0000001111000001",
"1101110111001011","1100010011101011","1100001100010010","1101101000110011",
"0000000001000000","0010011000110011","0011110100010010","0011110011101011",
"0010001111001011","1111110111000001","1101100011001111","1100001011110001",
"1100010100011000","1110000000110110","0000011000111111","0010101000101111",
"0011111000001100","0011100111100101","0001111011001000","1111011111000001",
"1101001111010011","1100000111110111","1100100000011110","1110010100111001",
"0000110000111110","0010111100101010","0011111100000110","0011011011100000",
"0001100011000101","1111000111000010","1100111111011000","1100000111111101",
"1100101100100011","1110101100111100","0001001000111101","0011001100100110",
"0100000000000000","0000100111000001","1100001111101110","1110010100111001",
"0011010100100011","0010101011010001","1101100011001111","1100101000100000",
"0001100000111011","0011111011110001","1111101011000001","1100000111111101",
"1111010000111110","0011110000010101","0001111011001000","1100110111011010",
"1101001100101101","0010011000110011","0011100011100010","1110101111000100",
"1100001000001100","0000001100111111","0011111100000110","0000111111000010",
"1100010111101000","1110000000110110","0011000100101000","0010111111010110",
"1101110111001011","1100011100011011","0001001000111101","0011111111110111",
"0000000011000000","1100000111110111","1110111000111101","0011100100011011",
"0010001111001011","1101000111010110","1100111100101000","0010000000110110",
"0011101111101000","1111000111000010","1100000100000110","1111110100111111",
"0011111000001100","0001010111000100","1100100011100010","1101101000110011",
"0010110100101101","0011001111011010","1110001011001000","1100010000010101",
"0000110000111110","0011111111111101","0000011011000001","1100001011110001",
"1110100000111011","0011011000100000","0010100011001111","1101011011010001",
"1100101100100011","0001101100111001","0011110111101110","1111011111000001",
"1100000000000000","1111011100111111","0011110100010010","0001101111000111",
"1100101111011101","1101011000101111","0010100000110001","0011011011100000",
"1110100011000101","1100001000001111","0000011000111111","0011111100000011",
"0000110011000010","1100010011101011","1110001000111000","0011001100100110",
"0010110111010011","1101101011001101","1100100000011110","0001010100111100",
"0011111011110100","1111110111000001","1100000111111010","1111000100111110",
"0011101100011000","0010000011001010","1100111111011000","1101000100101010",
"0010001100110101","0011100111100101","1110111011000011","1100000100001001",
"0000000001000000","0011111100001001","0001001011000011","1100011111100101",
"1101110100110101","0010111100101010","0011000111011000","1110000011001010",
"1100010100011000","0000111100111110","0011111111111010","0000001111000001",
"1100001011110100","1110101100111100","0011100000011110","0010011011001101",
"1101001111010011","1100110100100110","0001111000111000","0011110011101011",
"1111010011000010","1100000100000011","1111101000111111","0011111000001111",
"0001100011000101","1100101011100000","1101100000110001","0010101000101111",
"0011010111011101","1110010111000111","1100001100010010","0000100100111111",
"0100000000000000","1101101011001101","1110111000111101","0011110011101011",
"1100101111011101","0000001100111111","0011000111011000","1100001011110001",
"0001100000111011","0010000011001010","1100000100000110","0010101000101111",
"0000110011000010","1100011100011011","0011100000011110","1111011111000001",
"1101001100101101","0011111100001001","1110001011001000","1110010100111001",
"0011111011110100","1101000111010110","1111101000111111","0011011011100000",
"1100010111101000","0000111100111110","0010100011001111","1100000111111101",
"0010001100110101","0001010111000100","1100001100010010","0011001100100110",
"0000000011000000","1100110100100110","0011110100010010","1110101111000100",
"1101110100110101","0011111111111101","1101100011001111","1111000100111110",
"0011101111101000","1100101011100000","0000011000111111","0010111111010110",
"1100001011110100","0001101100111001","0001111011001000","1100000100001001",
"0010110100101101","0000100111000001","1100100000011110","0011100100011011",
"1111010011000010","1101011000101111","0011111100000110","1110000011001010",
"1110100000111011","0011111011110001","1100111111011000","1111110100111111",
"0011010111011101","1100010011101011","0001001000111101","0010011011001101",
"1100000000000000","0010011000110011","0001001011000011","1100010000010101",
"0011010100100011","1111110111000001","1100111100101000","0011111000001111",
"1110100011000101","1110000000110110","0011111111111010","1101011011010001",
"1111010000111110","0011100111100101","1100100011100010","0000100100111111",
"0010110111010011","1100000111110111","0001111000111000","0001101111000111",
"1100001000001100","0010111100101010","0000011011000001","1100101000100000",
"0011101100011000","1111000111000010","1101100000110001","0011111100000011",
"1101110111001011","1110101100111100","0011110111101110","1100110111011010",
"0000000001000000","0011001111011010","1100001111101110","0001010100111100",
"0010001111001011","1100000100000011","0010100000110001","0000111111000010",
"1100010100011000","0011011000100000","1111101011000001","1101000100101010",
"0011111000001100","1110010111000111","1110001000111000","0011111111110111",
"1101001111010011","1111011100111111","0011100011100010","1100011111100101",
"0000110000111110","0010101011010001","1100000111111010","0010000000110110",
"0001100011000101","1100001000001111","0011000100101000","0000001111000001",
"1100101100100011","0011110000010101","1110111011000011","1101101000110011",
"0100000000000000","1100000111110111","0011110100010010","1100011111100101",
"0011010100100011","1101000111010110","0010100000110001","1110000011001010",
"0001100000111011","1111000111000010","0000011000111111","0000001111000001",
"1111010000111110","0001010111000100","1110001000111000","0010011011001101",
"1101001100101101","0011001111011010","1100100000011110","0011110011101011",
"1100001000001100","0011111111111101","1100000111111010","0011111000001111",
"1100010111101000","0011011000100000","1100111111011000","0010101000101111",
"1101110111001011","0001101100111001","1110111011000011","0000100100111111",
"0000000011000000","1111011100111111","0001001011000011","1110010100111001",
"0010001111001011","1101011000101111","0011000111011000","1100101000100000",
"0011101111101000","1100001000001111","0011111111111010","1100000111111101",
"0011111000001100","1100010011101011","0011100000011110","1100110111011010",
"0010110100101101","1101101011001101","0001111000111000","1110101111000100",
"0000110000111110","1111110111000001","1111101000111111","0000111111000010",
"1110100000111011","0010000011001010","1101100000110001","0010111111010110",
"1100101100100011","0011100111100101","1100001100010010","0011111111110111",
"1100000000000000","0011111100001001","1100001111101110","0011100100011011",
"1100101111011101","0010111100101010","1101100011001111","0010000000110110",
"1110100011000101","0000111100111110","1111101011000001","1111110100111111",
"0000110011000010","1110101100111100","0001111011001000","1101101000110011",
"0010110111010011","1100110100100110","0011100011100010","1100010000010101",
"0011111011110100","1100000100000011","0011111100000110","1100001011110001",
"0011101100011000","1100101011100000","0011000100101000","1101011011010001",
"0010001100110101","1110010111000111","0001001000111101","1111011111000001",
"0000000001000000","0000100111000001","1110111000111101","0001101111000111",
"1101110100110101","0010101011010001","1100111100101000","0011011011100000",
"1100010100011000","0011111011110001","1100000100000110","0011111100000011",
"1100001011110100","0011110000010101","1100100011100010","0011001100100110",
"1101001111010011","0010011000110011","1110001011001000","0001010100111100",
"1111010011000010","0000001100111111","0000011011000001","1111000100111110",
"0001100011000101","1110000000110110","0010100011001111","1101000100101010",
"0011010111011101","1100011100011011","0011110111101110","1100000100001001"
),
("0100000000000000","0011000111011000","0000110011000010","1110001011001000",
"1100010111101000","1100001100010010","1101110100110101","0000011000111111",
"0010110100101101","0011111100000110","0011010111011101","0001001011000011",
"1110100011000101","1100100011100010","1100001000001100","1101100000110001",
"0000000001000000","0010100000110001","0011111000001100","0011100011100010",
"0001100011000101","1110111011000011","1100101111011101","1100000100000110",
"1101001100101101","1111101000111111","0010001100110101","0011110100010010",
"0011101111101000","0001111011001000","1111010011000010","1100111111011000",
"1100000000000000","1100111100101000","1111010000111110","0001111000111000",
"0011101100011000","0011110111101110","0010001111001011","1111101011000001",
"1101001111010011","1100000111111010","1100101100100011","1110111000111101",
"0001100000111011","0011100000011110","0011111011110100","0010100011001111",
"0000000011000000","1101100011001111","1100001011110100","1100100000011110",
"1110100000111011","0001001000111101","0011010100100011","0011111111111010",
"0010110111010011","0000011011000001","1101110111001011","1100001111101110",
"1100010100011000","1110001000111000","0000110000111110","0011000100101000",
"0100000000000000","0011000111011000","0000110011000010","1110001011001000",
"1100010111101000","1100001100010010","1101110100110101","0000011000111111",
"0010110100101101","0011111100000110","0011010111011101","0001001011000011",
"1110100011000101","1100100011100010","1100001000001100","1101100000110001",
"0000000001000000","0010100000110001","0011111000001100","0011100011100010",
"0001100011000101","1110111011000011","1100101111011101","1100000100000110",
"1101001100101101","1111101000111111","0010001100110101","0011110100010010",
"0011101111101000","0001111011001000","1111010011000010","1100111111011000",
"1100000000000000","1100111100101000","1111010000111110","0001111000111000",
"0011101100011000","0011110111101110","0010001111001011","1111101011000001",
"1101001111010011","1100000111111010","1100101100100011","1110111000111101",
"0001100000111011","0011100000011110","0011111011110100","0010100011001111",
"0000000011000000","1101100011001111","1100001011110100","1100100000011110",
"1110100000111011","0001001000111101","0011010100100011","0011111111111010",
"0010110111010011","0000011011000001","1101110111001011","1100001111101110",
"1100010100011000","1110001000111000","0000110000111110","0011000100101000",
"0100000000000000","0000011011000001","1100001011110100","1110111000111101",
"0011101100011000","0001111011001000","1100101111011101","1101100000110001",
"0010110100101101","0011000111011000","1101110111001011","1100100000011110",
"0001100000111011","0011110111101110","1111010011000010","1100000100000110",
"0000000001000000","0011111100000110","0000110011000010","1100001111101110",
"1110100000111011","0011100000011110","0010001111001011","1100111111011000",
"1101001100101101","0010100000110001","0011010111011101","1110001011001000",
"1100010100011000","0001001000111101","0011111011110100","1111101011000001",
"1100000000000000","1111101000111111","0011111000001100","0001001011000011",
"1100010111101000","1110001000111000","0011010100100011","0010100011001111",
"1101001111010011","1100111100101000","0010001100110101","0011100011100010",
"1110100011000101","1100001100010010","0000110000111110","0011111111111010",
"0000000011000000","1100000111111010","1111010000111110","0011110100010010",
"0001100011000101","1100100011100010","1101110100110101","0011000100101000",
"0010110111010011","1101100011001111","1100101100100011","0001111000111000",
"0011101111101000","1110111011000011","1100001000001100","0000011000111111",
"0100000000000000","0000011011000001","1100001011110100","1110111000111101",
"0011101100011000","0001111011001000","1100101111011101","1101100000110001",
"0010110100101101","0011000111011000","1101110111001011","1100100000011110",
"0001100000111011","0011110111101110","1111010011000010","1100000100000110",
"0000000001000000","0011111100000110","0000110011000010","1100001111101110",
"1110100000111011","0011100000011110","0010001111001011","1100111111011000",
"1101001100101101","0010100000110001","0011010111011101","1110001011001000",
"1100010100011000","0001001000111101","0011111011110100","1111101011000001",
"1100000000000000","1111101000111111","0011111000001100","0001001011000011",
"1100010111101000","1110001000111000","0011010100100011","0010100011001111",
"1101001111010011","1100111100101000","0010001100110101","0011100011100010",
"1110100011000101","1100001100010010","0000110000111110","0011111111111010",
"0000000011000000","1100000111111010","1111010000111110","0011110100010010",
"0001100011000101","1100100011100010","1101110100110101","0011000100101000",
"0010110111010011","1101100011001111","1100101100100011","0001111000111000",
"0011101111101000","1110111011000011","1100001000001100","0000011000111111",
"0100000000000000","1101100011001111","1111010000111110","0011100011100010",
"1100010111101000","0001001000111101","0010001111001011","1100000100000110",
"0010110100101101","0000011011000001","1100101100100011","0011110100010010",
"1110100011000101","1110001000111000","0011111011110100","1100111111011000",
"0000000001000000","0011000111011000","1100001011110100","0001111000111000",
"0001100011000101","1100001100010010","0011010100100011","1111101011000001",
"1101001100101101","0011111100000110","1101110111001011","1110111000111101",
"0011101111101000","1100100011100010","0000110000111110","0010100011001111",
"1100000000000000","0010100000110001","0000110011000010","1100100000011110",
"0011101100011000","1110111011000011","1101110100110101","0011111111111010",
"1101001111010011","1111101000111111","0011010111011101","1100001111101110",
"0001100000111011","0001111011001000","1100001000001100","0011000100101000",
"0000000011000000","1100111100101000","0011111000001100","1110001011001000",
"1110100000111011","0011110111101110","1100101111011101","0000011000111111",
"0010110111010011","1100000111111010","0010001100110101","0001001011000011",
"1100010100011000","0011100000011110","1111010011000010","1101100000110001",
"0100000000000000","1101100011001111","1111010000111110","0011100011100010",
"1100010111101000","0001001000111101","0010001111001011","1100000100000110",
"0010110100101101","0000011011000001","1100101100100011","0011110100010010",
"1110100011000101","1110001000111000","0011111011110100","1100111111011000",
"0000000001000000","0011000111011000","1100001011110100","0001111000111000",
"0001100011000101","1100001100010010","0011010100100011","1111101011000001",
"1101001100101101","0011111100000110","1101110111001011","1110111000111101",
"0011101111101000","1100100011100010","0000110000111110","0010100011001111",
"1100000000000000","0010100000110001","0000110011000010","1100100000011110",
"0011101100011000","1110111011000011","1101110100110101","0011111111111010",
"1101001111010011","1111101000111111","0011010111011101","1100001111101110",
"0001100000111011","0001111011001000","1100001000001100","0011000100101000",
"0000000011000000","1100111100101000","0011111000001100","1110001011001000",
"1110100000111011","0011110111101110","1100101111011101","0000011000111111",
"0010110111010011","1100000111111010","0010001100110101","0001001011000011",
"1100010100011000","0011100000011110","1111010011000010","1101100000110001",
"0100000000000000","1100000111111010","0011111000001100","1100001111101110",
"0011101100011000","1100100011100010","0011010100100011","1100111111011000",
"0010110100101101","1101100011001111","0010001100110101","1110001011001000",
"0001100000111011","1110111011000011","0000110000111110","1111101011000001",
"0000000001000000","0000011011000001","1111010000111110","0001001011000011",
"1110100000111011","0001111011001000","1101110100110101","0010100011001111",
"1101001100101101","0011000111011000","1100101100100011","0011100011100010",
"1100010100011000","0011110111101110","1100001000001100","0011111111111010",
"1100000000000000","0011111100000110","1100001011110100","0011110100010010",
"1100010111101000","0011100000011110","1100101111011101","0011000100101000",
"1101001111010011","0010100000110001","1101110111001011","0001111000111000",
"1110100011000101","0001001000111101","1111010011000010","0000011000111111",
"0000000011000000","1111101000111111","0000110011000010","1110111000111101",
"0001100011000101","1110001000111000","0010001111001011","1101100000110001",
"0010110111010011","1100111100101000","0011010111011101","1100100000011110",
"0011101111101000","1100001100010010","0011111011110100","1100000100000110",
"0100000000000000","1100000111111010","0011111000001100","1100001111101110",
"0011101100011000","1100100011100010","0011010100100011","1100111111011000",
"0010110100101101","1101100011001111","0010001100110101","1110001011001000",
"0001100000111011","1110111011000011","0000110000111110","1111101011000001",
"0000000001000000","0000011011000001","1111010000111110","0001001011000011",
"1110100000111011","0001111011001000","1101110100110101","0010100011001111",
"1101001100101101","0011000111011000","1100101100100011","0011100011100010",
"1100010100011000","0011110111101110","1100001000001100","0011111111111010",
"1100000000000000","0011111100000110","1100001011110100","0011110100010010",
"1100010111101000","0011100000011110","1100101111011101","0011000100101000",
"1101001111010011","0010100000110001","1101110111001011","0001111000111000",
"1110100011000101","0001001000111101","1111010011000010","0000011000111111",
"0000000011000000","1111101000111111","0000110011000010","1110111000111101",
"0001100011000101","1110001000111000","0010001111001011","1101100000110001",
"0010110111010011","1100111100101000","0011010111011101","1100100000011110",
"0011101111101000","1100001100010010","0011111011110100","1100000100000110"
),
("0100000000000000","0010111111010110","0000011011000001","1101101011001101",
"1100001011110100","1100101000100000","1110111000111101","0001101100111001",
"0011101100011000","0011110011101011","0001111011001000","1111000111000010",
"1100101111011101","1100000100001001","1101100000110001","0000001100111111",
"0010110100101101","0011111100000011","0011000111011000","0000100111000001",
"1101110111001011","1100001011110001","1100100000011110","1110101100111100",
"0001100000111011","0011100100011011","0011110111101110","0010000011001010",
"1111010011000010","1100110111011010","1100000100000110","1101011000101111",
"0000000001000000","0010101000101111","0011111100000110","0011001111011010",
"0000110011000010","1110000011001010","1100001111101110","1100011100011011",
"1110100000111011","0001010100111100","0011100000011110","0011111011110001",
"0010001111001011","1111011111000001","1100111111011000","1100000100000011",
"1101001100101101","1111110100111111","0010100000110001","0011111100001001",
"0011010111011101","0000111111000010","1110001011001000","1100010011101011",
"1100010100011000","1110010100111001","0001001000111101","0011011000100000",
"0011111011110100","0010011011001101","1111101011000001","1101000111010110",
"1100000000000000","1101000100101010","1111101000111111","0010011000110011",
"0011111000001100","0011011011100000","0001001011000011","1110010111000111",
"1100010111101000","1100010000010101","1110001000111000","0000111100111110",
"0011010100100011","0011111111110111","0010100011001111","1111110111000001",
"1101001111010011","1100000111111101","1100111100101000","1111011100111111",
"0010001100110101","0011111000001111","0011100011100010","0001010111000100",
"1110100011000101","1100011111100101","1100001100010010","1110000000110110",
"0000110000111110","0011001100100110","0011111111111010","0010101011010001",
"0000000011000000","1101011011010001","1100000111111010","1100110100100110",
"1111010000111110","0010000000110110","0011110100010010","0011100111100101",
"0001100011000101","1110101111000100","1100100011100010","1100001000001111",
"1101110100110101","0000100100111111","0011000100101000","0011111111111101",
"0010110111010011","0000001111000001","1101100011001111","1100000111110111",
"1100101100100011","1111000100111110","0001111000111000","0011110000010101",
"0011101111101000","0001101111000111","1110111011000011","1100101011100000",
"1100001000001100","1101101000110011","0000011000111111","0010111100101010",
"0100000000000000","0000001111000001","1100000111111010","1111011100111111",
"0011111000001100","0000111111000010","1100001111101110","1110101100111100",
"0011101100011000","0001101111000111","1100100011100010","1110000000110110",
"0011010100100011","0010011011001101","1100111111011000","1101011000101111",
"0010110100101101","0010111111010110","1101100011001111","1100110100100110",
"0010001100110101","0011011011100000","1110001011001000","1100011100011011",
"0001100000111011","0011110011101011","1110111011000011","1100001000001111",
"0000110000111110","0011111111110111","1111101011000001","1100000100000011",
"0000000001000000","0011111100000011","0000011011000001","1100000111110111",
"1111010000111110","0011111000001111","0001001011000011","1100010011101011",
"1110100000111011","0011100100011011","0001111011001000","1100101011100000",
"1101110100110101","0011001100100110","0010100011001111","1101000111010110",
"1101001100101101","0010101000101111","0011000111011000","1101101011001101",
"1100101100100011","0010000000110110","0011100011100010","1110010111000111",
"1100010100011000","0001010100111100","0011110111101110","1111000111000010",
"1100001000001100","0000100100111111","0011111111111010","1111110111000001",
"1100000000000000","1111110100111111","0011111100000110","0000100111000001",
"1100001011110100","1111000100111110","0011110100010010","0001010111000100",
"1100010111101000","1110010100111001","0011100000011110","0010000011001010",
"1100101111011101","1101101000110011","0011000100101000","0010101011010001",
"1101001111010011","1101000100101010","0010100000110001","0011001111011010",
"1101110111001011","1100101000100000","0001111000111000","0011100111100101",
"1110100011000101","1100010000010101","0001001000111101","0011111011110001",
"1111010011000010","1100000100001001","0000011000111111","0011111111111101",
"0000000011000000","1100000111111101","1111101000111111","0011111100001001",
"0000110011000010","1100001011110001","1110111000111101","0011110000010101",
"0001100011000101","1100011111100101","1110001000111000","0011011000100000",
"0010001111001011","1100110111011010","1101100000110001","0010111100101010",
"0010110111010011","1101011011010001","1100111100101000","0010011000110011",
"0011010111011101","1110000011001010","1100100000011110","0001101100111001",
"0011101111101000","1110101111000100","1100001100010010","0000111100111110",
"0011111011110100","1111011111000001","1100000100000110","0000001100111111",
"0100000000000000","1101011011010001","1111101000111111","0011001111011010",
"1100001011110100","0010000000110110","0001001011000011","1100011100011011",
"0011101100011000","1110101111000100","1110001000111000","0011111011110001",
"1100101111011101","0000100100111111","0010100011001111","1100000100000011",
"0010110100101101","0000001111000001","1100111100101000","0011111100001001",
"1101110111001011","1111000100111110","0011100011100010","1100010011101011",
"0001100000111011","0001101111000111","1100001100010010","0011011000100000",
"1111010011000010","1101101000110011","0011111111111010","1101000111010110",
"0000000001000000","0010111111010110","1100000111111010","0010011000110011",
"0000110011000010","1100101000100000","0011110100010010","1110010111000111",
"1110100000111011","0011110011101011","1100100011100010","0000111100111110",
"0010001111001011","1100000100001001","0011000100101000","1111110111000001",
"1101001100101101","0011111100000011","1101100011001111","1111011100111111",
"0011010111011101","1100001011110001","0001111000111000","0001010111000100",
"1100010100011000","0011100100011011","1110111011000011","1110000000110110",
"0011111011110100","1100110111011010","0000011000111111","0010101011010001",
"1100000000000000","0010101000101111","0000011011000001","1100110100100110",
"0011111000001100","1110000011001010","1110111000111101","0011100111100101",
"1100010111101000","0001010100111100","0001111011001000","1100001000001111",
"0011010100100011","1111011111000001","1101100000110001","0011111111111101",
"1101001111010011","1111110100111111","0011000111011000","1100000111110111",
"0010001100110101","0000111111000010","1100100000011110","0011110000010101",
"1110100011000101","1110010100111001","0011110111101110","1100101011100000",
"0000110000111110","0010011011001101","1100000100000110","0010111100101010",
"0000000011000000","1101000100101010","0011111100000110","1101101011001101",
"1111010000111110","0011011011100000","1100001111101110","0001101100111001",
"0001100011000101","1100010000010101","0011100000011110","1111000111000010",
"1101110100110101","0011111111110111","1100111111011000","0000001100111111",
"0010110111010011","1100000111111101","0010100000110001","0000100111000001",
"1100101100100011","0011111000001111","1110001011001000","1110101100111100",
"0011101111101000","1100011111100101","0001001000111101","0010000011001010",
"1100001000001100","0011001100100110","1111101011000001","1101011000101111",
"0100000000000000","1100000111111101","0011111100000110","1100000111110111",
"0011111000001100","1100001011110001","0011110100010010","1100010011101011",
"0011101100011000","1100011111100101","0011100000011110","1100101011100000",
"0011010100100011","1100110111011010","0011000100101000","1101000111010110",
"0010110100101101","1101011011010001","0010100000110001","1101101011001101",
"0010001100110101","1110000011001010","0001111000111000","1110010111000111",
"0001100000111011","1110101111000100","0001001000111101","1111000111000010",
"0000110000111110","1111011111000001","0000011000111111","1111110111000001",
"0000000001000000","0000001111000001","1111101000111111","0000100111000001",
"1111010000111110","0000111111000010","1110111000111101","0001010111000100",
"1110100000111011","0001101111000111","1110001000111000","0010000011001010",
"1101110100110101","0010011011001101","1101100000110001","0010101011010001",
"1101001100101101","0010111111010110","1100111100101000","0011001111011010",
"1100101100100011","0011011011100000","1100100000011110","0011100111100101",
"1100010100011000","0011110011101011","1100001100010010","0011111011110001",
"1100001000001100","0011111111110111","1100000100000110","0011111111111101",
"1100000000000000","0011111100000011","1100000111111010","0011111100001001",
"1100001011110100","0011111000001111","1100001111101110","0011110000010101",
"1100010111101000","0011100100011011","1100100011100010","0011011000100000",
"1100101111011101","0011001100100110","1100111111011000","0010111100101010",
"1101001111010011","0010101000101111","1101100011001111","0010011000110011",
"1101110111001011","0010000000110110","1110001011001000","0001101100111001",
"1110100011000101","0001010100111100","1110111011000011","0000111100111110",
"1111010011000010","0000100100111111","1111101011000001","0000001100111111",
"0000000011000000","1111110100111111","0000011011000001","1111011100111111",
"0000110011000010","1111000100111110","0001001011000011","1110101100111100",
"0001100011000101","1110010100111001","0001111011001000","1110000000110110",
"0010001111001011","1101101000110011","0010100011001111","1101011000101111",
"0010110111010011","1101000100101010","0011000111011000","1100110100100110",
"0011010111011101","1100101000100000","0011100011100010","1100011100011011",
"0011101111101000","1100010000010101","0011110111101110","1100001000001111",
"0011111011110100","1100000100001001","0011111111111010","1100000100000011"
));
end twiddles;
