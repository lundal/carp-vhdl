-------------------------------------------------------------------------------
-- Title      : Toplevel
-- Project    : Cellular Automata Research Platform
-------------------------------------------------------------------------------
-- File       : toplevel.vhd
-- Author     : Per Thomas Lundal <perthomas@gmail.com>
-- Company    : NTNU
-- Last update: 2015-01-20
-- Platform   : Spartan-6
-------------------------------------------------------------------------------
-- Description: Connects all main components
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author    Description
-- 2015-01-20  1.0      lundal    Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.functions.all;
use work.types.all;

entity toplevel is
  generic (
    tx_buffer_address_bits   : positive := 10; -- PCIe packet length field is 10 bits
    rx_buffer_address_bits   : positive := 10;
    reverse_payload_endian   : boolean  := true; -- Required for x86 systems
    program_counter_bits     : positive := 8;
    matrix_width             : positive := 8;
    matrix_height            : positive := 8;
    matrix_depth             : positive := 8;
    matrix_wrap              : boolean  := true;
    cell_type_bits           : positive := 8;
    cell_state_bits          : positive := 1; -- Must be 1 due to implementation of CA
    jump_counters            : positive := 4;
    jump_counter_bits        : positive := 16;
    instruction_bits         : positive := 256; -- Must be 256 due to implementation of fetch_communication
    lut_configuration_bits   : positive := 8; -- Should optimally be 2 for 2D and 8 for 3D
    rule_vector_amount       : positive := 64;
    rule_amount              : positive := 256;
    rules_tested_in_parallel : positive := 4;
    live_count_buffer_size   : positive := 256;
    fitness_buffer_size      : positive := 256
  );
  port (
    pcie_tx_p : out std_logic;
    pcie_tx_n : out std_logic;
    pcie_rx_p : in  std_logic;
    pcie_rx_n : in  std_logic;

    clock_p : in  std_logic;
    clock_n : in  std_logic;
    reset_n : in  std_logic;

    leds : out std_logic_vector(3 downto 0)
  );
end toplevel;

architecture rtl of toplevel is

  -- Calculate amount of cells that fits in one write instruction
  constant cell_type_write_width  : positive := min(matrix_width, (instruction_bits-32)/cell_type_bits);
  constant cell_state_write_width : positive := min(matrix_width, (instruction_bits-32)/cell_state_bits);

  -- Inferred constants
  constant live_count_buffer_bits : positive := bits(matrix_depth*matrix_height*matrix_width) + 1; -- From cellular automata
  constant send_buffer_size       : positive := 2**tx_buffer_address_bits;

  -- General
  signal clock : std_logic;
  signal reset : std_logic;

  -- Pipeline control
  signal run                      : std_logic;
  signal done_fetch               : std_logic;
  signal done_information_sender  : std_logic;
  signal done_cell_writer_reader  : std_logic;
  signal done_cellular_automata   : std_logic;
  signal done_development         : std_logic;
  signal done_rule_vector_reader  : std_logic;
  signal done_rule_numbers_reader : std_logic;
  signal done_fitness_sender      : std_logic;

  -- Communication
  signal tx_buffer_data  : std_logic_vector(31 downto 0);
  signal tx_buffer_count : std_logic_vector(tx_buffer_address_bits - 1 downto 0);
  signal tx_buffer_write : std_logic;

  signal rx_buffer_data  : std_logic_vector(31 downto 0);
  signal rx_buffer_count : std_logic_vector(rx_buffer_address_bits - 1 downto 0);
  signal rx_buffer_read  : std_logic;

  -- Decode
  signal decode_from_fetch_instruction : std_logic_vector(instruction_bits - 1 downto 0);

  signal decode_to_information_sender_operation : information_sender_operation_type;

  signal decode_to_cell_writer_reader_operation : cell_writer_reader_operation_type;
  signal decode_to_cell_writer_reader_address_z : std_logic_vector(bits(matrix_depth) - 1 downto 0);
  signal decode_to_cell_writer_reader_address_y : std_logic_vector(bits(matrix_height) - 1 downto 0);
  signal decode_to_cell_writer_reader_address_x : std_logic_vector(bits(matrix_width) - 1 downto 0);
  signal decode_to_cell_writer_reader_state     : std_logic_vector(cell_state_bits - 1 downto 0);
  signal decode_to_cell_writer_reader_states    : std_logic_vector(cell_state_write_width*cell_state_bits - 1 downto 0);
  signal decode_to_cell_writer_reader_type      : std_logic_vector(cell_type_bits - 1 downto 0);
  signal decode_to_cell_writer_reader_types     : std_logic_vector(cell_type_write_width*cell_type_bits - 1 downto 0);

  signal decode_to_cellular_automata_operation  : cellular_automata_operation_type;
  signal decode_to_cellular_automata_step_count : std_logic_vector(15 downto 0);

  signal decode_to_development_operation    : development_operation_type;
  signal decode_to_development_rules_active : std_logic_vector(bits(rule_amount) - 1 downto 0);

  signal decode_to_lut_writer_operation : lut_writer_operation_type;
  signal decode_to_lut_writer_address   : std_logic_vector(cell_type_bits - 1 downto 0);
  signal decode_to_lut_writer_data      : std_logic_vector(2**if_else(matrix_depth = 1, 5, 7) - 1 downto 0);

  signal decode_to_rule_writer_operation : rule_writer_operation_type;
  signal decode_to_rule_writer_address   : std_logic_vector(bits(rule_amount) - 1 downto 0);
  signal decode_to_rule_writer_data      : std_logic_vector((cell_type_bits + 1 + cell_state_bits + 1) * if_else(matrix_depth = 1, 6, 8) - 1 downto 0);

  signal decode_to_rule_vector_reader_operation : rule_vector_reader_operation_type;
  signal decode_to_rule_vector_reader_count     : std_logic_vector(bits(rule_vector_amount) - 1 downto 0);

  signal decode_to_rule_numbers_reader_operation : rule_numbers_reader_operation_type;

  signal decode_to_fitness_sender_operation : fitness_sender_operation_type;

  signal decode_to_buffers_reset          : std_logic;
  signal decode_to_cell_buffer_swap       : std_logic;
  signal decode_to_cell_buffer_mux_select : cell_buffer_mux_select_type;
  signal decode_to_send_buffer_mux_select : send_buffer_mux_select_type;

  -- Information Sender
  signal information_sender_to_send_mux_data    : std_logic_vector(31 downto 0);
  signal information_sender_from_send_mux_count : std_logic_vector(tx_buffer_address_bits - 1 downto 0);
  signal information_sender_to_send_mux_write   : std_logic;

  -- Cell Writer Reader
  signal cell_writer_reader_to_mux_address_z    : std_logic_vector(bits(matrix_depth) - 1 downto 0);
  signal cell_writer_reader_to_mux_address_y    : std_logic_vector(bits(matrix_height) - 1 downto 0);
  signal cell_writer_reader_to_mux_types_write  : std_logic;
  signal cell_writer_reader_to_mux_types        : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal cell_writer_reader_from_mux_types      : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal cell_writer_reader_to_mux_states_write : std_logic;
  signal cell_writer_reader_to_mux_states       : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);
  signal cell_writer_reader_from_mux_states     : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);

  signal cell_writer_reader_to_send_mux_data    : std_logic_vector(31 downto 0);
  signal cell_writer_reader_from_send_mux_count : std_logic_vector(tx_buffer_address_bits - 1 downto 0);
  signal cell_writer_reader_to_send_mux_write   : std_logic;

  -- Cellular Automata
  signal cellular_automata_to_mux_address_z    : std_logic_vector(bits(matrix_depth) - 1 downto 0);
  signal cellular_automata_to_mux_address_y    : std_logic_vector(bits(matrix_height) - 1 downto 0);
  signal cellular_automata_to_mux_types_write  : std_logic;
  signal cellular_automata_to_mux_types        : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal cellular_automata_from_mux_types      : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal cellular_automata_to_mux_states_write : std_logic;
  signal cellular_automata_to_mux_states       : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);
  signal cellular_automata_from_mux_states     : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);

  -- Development
  signal development_to_mux_a_address_z    : std_logic_vector(bits(matrix_depth) - 1 downto 0);
  signal development_to_mux_a_address_y    : std_logic_vector(bits(matrix_height) - 1 downto 0);
  signal development_to_mux_a_types_write  : std_logic;
  signal development_to_mux_a_types        : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal development_from_mux_a_types      : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal development_to_mux_a_states_write : std_logic;
  signal development_to_mux_a_states       : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);
  signal development_from_mux_a_states     : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);

  signal development_to_mux_b_address_z    : std_logic_vector(bits(matrix_depth) - 1 downto 0);
  signal development_to_mux_b_address_y    : std_logic_vector(bits(matrix_height) - 1 downto 0);
  signal development_to_mux_b_types_write  : std_logic;
  signal development_to_mux_b_types        : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal development_from_mux_b_types      : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal development_to_mux_b_states_write : std_logic;
  signal development_to_mux_b_states       : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);
  signal development_from_mux_b_states     : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);

  -- Cell buffer
  signal cell_buffer_from_mux_a_address_z    : std_logic_vector(bits(matrix_depth) - 1 downto 0);
  signal cell_buffer_from_mux_a_address_y    : std_logic_vector(bits(matrix_height) - 1 downto 0);
  signal cell_buffer_from_mux_a_types_write  : std_logic;
  signal cell_buffer_from_mux_a_types        : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal cell_buffer_to_mux_a_types          : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal cell_buffer_from_mux_a_states_write : std_logic;
  signal cell_buffer_from_mux_a_states       : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);
  signal cell_buffer_to_mux_a_states         : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);

  signal cell_buffer_from_mux_b_address_z    : std_logic_vector(bits(matrix_depth) - 1 downto 0);
  signal cell_buffer_from_mux_b_address_y    : std_logic_vector(bits(matrix_height) - 1 downto 0);
  signal cell_buffer_from_mux_b_types_write  : std_logic;
  signal cell_buffer_from_mux_b_types        : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal cell_buffer_to_mux_b_types          : std_logic_vector(matrix_width*cell_type_bits - 1 downto 0);
  signal cell_buffer_from_mux_b_states_write : std_logic;
  signal cell_buffer_from_mux_b_states       : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);
  signal cell_buffer_to_mux_b_states         : std_logic_vector(matrix_width*cell_state_bits - 1 downto 0);

  -- LUT writer
  signal lut_writer_to_cellular_automata_write   : std_logic;
  signal lut_writer_to_cellular_automata_address : std_logic_vector(cell_type_bits - 1 downto 0);
  signal lut_writer_to_cellular_automata_data    : std_logic_vector(2**if_else(matrix_depth = 1, 5, 7) - 1 downto 0);

  -- Rule writer
  signal rule_writer_to_development_write   : std_logic;
  signal rule_writer_to_development_address : std_logic_vector(bits(rule_amount) - 1 downto 0);
  signal rule_writer_to_development_data    : std_logic_vector((cell_type_bits + 1 + cell_state_bits + 1) * if_else(matrix_depth = 1, 6, 8) - 1 downto 0);

  -- Rule vector reader
  signal rule_vector_reader_from_development_data  : std_logic_vector(rule_amount - 1 downto 0);
  signal rule_vector_reader_from_development_count : std_logic_vector(bits(rule_vector_amount) - 1 downto 0);
  signal rule_vector_reader_to_development_read    : std_logic;

  signal rule_vector_reader_to_send_mux_data    : std_logic_vector(31 downto 0);
  signal rule_vector_reader_from_send_mux_count : std_logic_vector(tx_buffer_address_bits - 1 downto 0);
  signal rule_vector_reader_to_send_mux_write   : std_logic;

  -- Rule numbers reader
  signal rule_numbers_reader_to_development_address_z : std_logic_vector(bits(matrix_depth) - 1 downto 0);
  signal rule_numbers_reader_to_development_address_y : std_logic_vector(bits(matrix_height) - 1 downto 0);
  signal rule_numbers_reader_from_development_data    : std_logic_vector(matrix_width * bits(rule_amount) - 1 downto 0);

  signal rule_numbers_reader_to_send_mux_data    : std_logic_vector(31 downto 0);
  signal rule_numbers_reader_from_send_mux_count : std_logic_vector(tx_buffer_address_bits - 1 downto 0);
  signal rule_numbers_reader_to_send_mux_write   : std_logic;

  -- Fitness
  signal fitness_to_live_count_buffer_read    : std_logic;
  signal fitness_from_live_count_buffer_data  : std_logic_vector(live_count_buffer_bits - 1 downto 0);
  signal fitness_from_live_count_buffer_count : std_logic_vector(bits(live_count_buffer_size) - 1 downto 0);

  signal fitness_to_buffer_write : std_logic;
  signal fitness_to_buffer_data  : std_logic_vector(32 - 1 downto 0);

  signal fitness_identifier    : std_logic_vector(8 - 1 downto 0);
  signal fitness_words_per_run : std_logic_vector(8 - 1 downto 0);
  signal fitness_parameters    : std_logic_vector(16 - 1 downto 0);

  -- Fitness buffer
  signal fitness_buffer_count : std_logic_vector(bits(fitness_buffer_size) - 1 downto 0);

  -- Fitness sender
  signal fitness_sender_to_send_mux_write   : std_logic;
  signal fitness_sender_to_send_mux_data    : std_logic_vector(32 - 1 downto 0);
  signal fitness_sender_from_send_mux_count : std_logic_vector(bits(send_buffer_size) - 1 downto 0);

  signal fitness_sender_to_buffer_read    : std_logic;
  signal fitness_sender_from_buffer_data  : std_logic_vector(32 - 1 downto 0);

begin

  leds <= "0101";

  run <= done_fetch
     and done_information_sender
     and done_cell_writer_reader
     and done_cellular_automata
     and done_development
     and done_rule_vector_reader
     and done_rule_numbers_reader
     and done_fitness_sender;

  -----------------------------------------------------------------------------

  communication : entity work.communication
  generic map (
    tx_buffer_address_bits => tx_buffer_address_bits,
    rx_buffer_address_bits => rx_buffer_address_bits,
    reverse_payload_endian => reverse_payload_endian
  )
  port map (
    pcie_tx_p => pcie_tx_p,
    pcie_tx_n => pcie_tx_n,
    pcie_rx_p => pcie_rx_p,
    pcie_rx_n => pcie_rx_n,

    clock_p => clock_p,
    clock_n => clock_n,
    reset_n => reset_n,

    tx_buffer_in    => tx_buffer_data,
    tx_buffer_count => tx_buffer_count,
    tx_buffer_write => tx_buffer_write,

    rx_buffer_out   => rx_buffer_data,
    rx_buffer_count => rx_buffer_count,
    rx_buffer_read  => rx_buffer_read,

    clock => clock,
    reset => reset
  );

  fetch : entity work.fetch
  generic map (
    buffer_address_bits  => rx_buffer_address_bits,
    jump_counters        => jump_counters,
    jump_counter_bits    => jump_counter_bits,
    program_counter_bits => program_counter_bits,
    instruction_bits     => instruction_bits
  )
  port map (
    buffer_data  => rx_buffer_data,
    buffer_count => rx_buffer_count,
    buffer_read  => rx_buffer_read,

    instruction => decode_from_fetch_instruction,

    run  => run,
    done => done_fetch,

    clock => clock
  );

  decode : entity work.decode
  generic map (
    matrix_width           => matrix_width,
    matrix_height          => matrix_height,
    matrix_depth           => matrix_depth,
    cell_type_bits         => cell_type_bits,
    cell_state_bits        => cell_state_bits,
    cell_type_write_width  => cell_type_write_width,
    cell_state_write_width => cell_state_write_width,
    instruction_bits       => instruction_bits,
    rule_amount            => rule_amount,
    rule_vector_amount     => rule_vector_amount
  )
  port map (
    instruction => decode_from_fetch_instruction,

    information_sender_operation => decode_to_information_sender_operation,

    cell_writer_reader_operation => decode_to_cell_writer_reader_operation,
    cell_writer_reader_address_z => decode_to_cell_writer_reader_address_z,
    cell_writer_reader_address_y => decode_to_cell_writer_reader_address_y,
    cell_writer_reader_address_x => decode_to_cell_writer_reader_address_x,
    cell_writer_reader_state     => decode_to_cell_writer_reader_state,
    cell_writer_reader_states    => decode_to_cell_writer_reader_states,
    cell_writer_reader_type      => decode_to_cell_writer_reader_type,
    cell_writer_reader_types     => decode_to_cell_writer_reader_types,

    cellular_automata_operation  => decode_to_cellular_automata_operation,
    cellular_automata_step_count => decode_to_cellular_automata_step_count,

    development_operation    => decode_to_development_operation,
    development_rules_active => decode_to_development_rules_active,

    lut_writer_operation => decode_to_lut_writer_operation,
    lut_writer_address   => decode_to_lut_writer_address,
    lut_writer_data      => decode_to_lut_writer_data,

    rule_writer_operation => decode_to_rule_writer_operation,
    rule_writer_address   => decode_to_rule_writer_address,
    rule_writer_data      => decode_to_rule_writer_data,

    rule_vector_reader_operation => decode_to_rule_vector_reader_operation,
    rule_vector_reader_count     => decode_to_rule_vector_reader_count,

    rule_numbers_reader_operation => decode_to_rule_numbers_reader_operation,

    fitness_sender_operation => decode_to_fitness_sender_operation,

    buffer_reset           => decode_to_buffers_reset,
    cell_buffer_swap       => decode_to_cell_buffer_swap,
    cell_buffer_mux_select => decode_to_cell_buffer_mux_select,
    send_buffer_mux_select => decode_to_send_buffer_mux_select,

    run  => run,

    clock => clock
  );

  information_sender : entity work.information_sender
  generic map (
    matrix_width             => matrix_width,
    matrix_height            => matrix_height,
    matrix_depth             => matrix_depth,
    matrix_wrap              => matrix_wrap,
    cell_type_bits           => cell_type_bits,
    cell_state_bits          => cell_state_bits,
    jump_counters            => jump_counters,
    jump_counter_bits        => jump_counter_bits,
    rule_amount              => rule_amount,
    send_buffer_address_bits => tx_buffer_address_bits
  )
  port map (
    send_buffer_data  => information_sender_to_send_mux_data,
    send_buffer_count => information_sender_from_send_mux_count,
    send_buffer_write => information_sender_to_send_mux_write,

    fitness_identifier    => fitness_identifier,
    fitness_words_per_run => fitness_words_per_run,
    fitness_parameters    => fitness_parameters,

    decode_operation => decode_to_information_sender_operation,

    run  => run,
    done => done_information_sender,

    clock => clock
  );

  cell_writer_reader : entity work.cell_writer_reader
  generic map (
    matrix_width             => matrix_width,
    matrix_height            => matrix_height,
    matrix_depth             => matrix_depth,
    cell_type_bits           => cell_type_bits,
    cell_state_bits          => cell_state_bits,
    cell_type_write_width    => cell_type_write_width,
    cell_state_write_width   => cell_state_write_width,
    send_buffer_address_bits => tx_buffer_address_bits
  )
  port map (
    buffer_address_z    => cell_writer_reader_to_mux_address_z,
    buffer_address_y    => cell_writer_reader_to_mux_address_y,
    buffer_types_write  => cell_writer_reader_to_mux_types_write,
    buffer_types_in     => cell_writer_reader_from_mux_types,
    buffer_types_out    => cell_writer_reader_to_mux_types,
    buffer_states_write => cell_writer_reader_to_mux_states_write,
    buffer_states_in    => cell_writer_reader_from_mux_states,
    buffer_states_out   => cell_writer_reader_to_mux_states,

    send_buffer_data  => cell_writer_reader_to_send_mux_data,
    send_buffer_count => cell_writer_reader_from_send_mux_count,
    send_buffer_write => cell_writer_reader_to_send_mux_write,

    decode_operation => decode_to_cell_writer_reader_operation,
    decode_address_z => decode_to_cell_writer_reader_address_z,
    decode_address_y => decode_to_cell_writer_reader_address_y,
    decode_address_x => decode_to_cell_writer_reader_address_x,
    decode_state     => decode_to_cell_writer_reader_state,
    decode_states    => decode_to_cell_writer_reader_states,
    decode_type      => decode_to_cell_writer_reader_type,
    decode_types     => decode_to_cell_writer_reader_types,

    run  => run,
    done => done_cell_writer_reader,

    clock => clock
  );

  cell_buffer_mux : entity work.cell_buffer_mux
  generic map (
    matrix_width    => matrix_width,
    matrix_height   => matrix_height,
    matrix_depth    => matrix_depth,
    cell_type_bits  => cell_type_bits,
    cell_state_bits => cell_state_bits
  )
  port map (
    writer_reader_address_z    => cell_writer_reader_to_mux_address_z,
    writer_reader_address_y    => cell_writer_reader_to_mux_address_y,
    writer_reader_types_write  => cell_writer_reader_to_mux_types_write,
    writer_reader_types_in     => cell_writer_reader_to_mux_types,
    writer_reader_types_out    => cell_writer_reader_from_mux_types,
    writer_reader_states_write => cell_writer_reader_to_mux_states_write,
    writer_reader_states_in    => cell_writer_reader_to_mux_states,
    writer_reader_states_out   => cell_writer_reader_from_mux_states,

    cellular_automata_address_z    => cellular_automata_to_mux_address_z,
    cellular_automata_address_y    => cellular_automata_to_mux_address_y,
    cellular_automata_types_write  => cellular_automata_to_mux_types_write,
    cellular_automata_types_in     => cellular_automata_to_mux_types,
    cellular_automata_types_out    => cellular_automata_from_mux_types,
    cellular_automata_states_write => cellular_automata_to_mux_states_write,
    cellular_automata_states_in    => cellular_automata_to_mux_states,
    cellular_automata_states_out   => cellular_automata_from_mux_states,

    development_a_address_z    => development_to_mux_a_address_z,
    development_a_address_y    => development_to_mux_a_address_y,
    development_a_types_write  => development_to_mux_a_types_write,
    development_a_types_in     => development_to_mux_a_types,
    development_a_types_out    => development_from_mux_a_types,
    development_a_states_write => development_to_mux_a_states_write,
    development_a_states_in    => development_to_mux_a_states,
    development_a_states_out   => development_from_mux_a_states,

    development_b_address_z    => development_to_mux_b_address_z,
    development_b_address_y    => development_to_mux_b_address_y,
    development_b_types_write  => development_to_mux_b_types_write,
    development_b_types_in     => development_to_mux_b_types,
    development_b_types_out    => development_from_mux_b_types,
    development_b_states_write => development_to_mux_b_states_write,
    development_b_states_in    => development_to_mux_b_states,
    development_b_states_out   => development_from_mux_b_states,

    buffer_a_address_z    => cell_buffer_from_mux_a_address_z,
    buffer_a_address_y    => cell_buffer_from_mux_a_address_y,
    buffer_a_types_write  => cell_buffer_from_mux_a_types_write,
    buffer_a_types_in     => cell_buffer_to_mux_a_types,
    buffer_a_types_out    => cell_buffer_from_mux_a_types,
    buffer_a_states_write => cell_buffer_from_mux_a_states_write,
    buffer_a_states_in    => cell_buffer_to_mux_a_states,
    buffer_a_states_out   => cell_buffer_from_mux_a_states,

    buffer_b_address_z    => cell_buffer_from_mux_b_address_z,
    buffer_b_address_y    => cell_buffer_from_mux_b_address_y,
    buffer_b_types_write  => cell_buffer_from_mux_b_types_write,
    buffer_b_types_in     => cell_buffer_to_mux_b_types,
    buffer_b_types_out    => cell_buffer_from_mux_b_types,
    buffer_b_states_write => cell_buffer_from_mux_b_states_write,
    buffer_b_states_in    => cell_buffer_to_mux_b_states,
    buffer_b_states_out   => cell_buffer_from_mux_b_states,

    source_select => decode_to_cell_buffer_mux_select,

    run => run,

    clock => clock
  );

  cell_buffer : entity work.cell_buffer
  generic map (
    matrix_width    => matrix_width,
    matrix_height   => matrix_height,
    matrix_depth    => matrix_depth,
    cell_type_bits  => cell_type_bits,
    cell_state_bits => cell_state_bits
  )
  port map (
    a_address_z    => cell_buffer_from_mux_a_address_z,
    a_address_y    => cell_buffer_from_mux_a_address_y,
    a_types_write  => cell_buffer_from_mux_a_types_write,
    a_types_in     => cell_buffer_from_mux_a_types,
    a_types_out    => cell_buffer_to_mux_a_types,
    a_states_write => cell_buffer_from_mux_a_states_write,
    a_states_in    => cell_buffer_from_mux_a_states,
    a_states_out   => cell_buffer_to_mux_a_states,

    b_address_z    => cell_buffer_from_mux_b_address_z,
    b_address_y    => cell_buffer_from_mux_b_address_y,
    b_types_write  => cell_buffer_from_mux_b_types_write,
    b_types_in     => cell_buffer_from_mux_b_types,
    b_types_out    => cell_buffer_to_mux_b_types,
    b_states_write => cell_buffer_from_mux_b_states_write,
    b_states_in    => cell_buffer_from_mux_b_states,
    b_states_out   => cell_buffer_to_mux_b_states,

    swap => decode_to_cell_buffer_swap,

    run => run,

    clock => clock
  );

  send_buffer_mux : entity work.send_buffer_mux
  generic map (
    send_buffer_address_bits => tx_buffer_address_bits
  )
  port map (
    cell_writer_reader_data  => cell_writer_reader_to_send_mux_data,
    cell_writer_reader_count => cell_writer_reader_from_send_mux_count,
    cell_writer_reader_write => cell_writer_reader_to_send_mux_write,

    information_sender_data  => information_sender_to_send_mux_data,
    information_sender_count => information_sender_from_send_mux_count,
    information_sender_write => information_sender_to_send_mux_write,

    rule_vector_reader_data  => rule_vector_reader_to_send_mux_data,
    rule_vector_reader_count => rule_vector_reader_from_send_mux_count,
    rule_vector_reader_write => rule_vector_reader_to_send_mux_write,

    rule_numbers_reader_data  => rule_numbers_reader_to_send_mux_data,
    rule_numbers_reader_count => rule_numbers_reader_from_send_mux_count,
    rule_numbers_reader_write => rule_numbers_reader_to_send_mux_write,

    fitness_sender_data  => fitness_sender_to_send_mux_data,
    fitness_sender_count => fitness_sender_from_send_mux_count,
    fitness_sender_write => fitness_sender_to_send_mux_write,

    send_buffer_data  => tx_buffer_data,
    send_buffer_count => tx_buffer_count,
    send_buffer_write => tx_buffer_write,

    source_select => decode_to_send_buffer_mux_select,

    run => run,

    clock => clock
  );

  cellular_automata : entity work.cellular_automata
  generic map (
    matrix_width           => matrix_width,
    matrix_height          => matrix_height,
    matrix_depth           => matrix_depth,
    matrix_wrap            => matrix_wrap,
    cell_type_bits         => cell_type_bits,
    cell_state_bits        => cell_state_bits,
    lut_configuration_bits => lut_configuration_bits,
    live_count_buffer_size => live_count_buffer_size
  )
  port map (
    buffer_address_z    => cellular_automata_to_mux_address_z,
    buffer_address_y    => cellular_automata_to_mux_address_y,
    buffer_types_write  => cellular_automata_to_mux_types_write,
    buffer_types_in     => cellular_automata_from_mux_types,
    buffer_types_out    => cellular_automata_to_mux_types,
    buffer_states_write => cellular_automata_to_mux_states_write,
    buffer_states_in    => cellular_automata_from_mux_states,
    buffer_states_out   => cellular_automata_to_mux_states,

    lut_storage_write   => lut_writer_to_cellular_automata_write,
    lut_storage_address => lut_writer_to_cellular_automata_address,
    lut_storage_data    => lut_writer_to_cellular_automata_data,

    live_count_read  => fitness_to_live_count_buffer_read,
    live_count_data  => fitness_from_live_count_buffer_data,
    live_count_count => fitness_from_live_count_buffer_count,
    live_count_reset => decode_to_buffers_reset,

    decode_operation  => decode_to_cellular_automata_operation,
    decode_step_count => decode_to_cellular_automata_step_count,

    run  => run,
    done => done_cellular_automata,

    clock => clock
  );

  lut_writer : entity work.lut_writer
  generic map (
    cell_type_bits => cell_type_bits,
    neighborhood_bits => if_else(matrix_depth = 1, 5, 7)
  )
  port map (
    lut_storage_write   => lut_writer_to_cellular_automata_write,
    lut_storage_address => lut_writer_to_cellular_automata_address,
    lut_storage_data    => lut_writer_to_cellular_automata_data,

    decode_operation => decode_to_lut_writer_operation,
    decode_address   => decode_to_lut_writer_address,
    decode_data      => decode_to_lut_writer_data,

    run => run,

    clock => clock
  );

  rule_writer : entity work.rule_writer
  generic map (
    cell_state_bits   => cell_state_bits,
    cell_type_bits    => cell_type_bits,
    neighborhood_size => if_else(matrix_depth = 1, 5, 7),
    rule_amount       => rule_amount
  )
  port map (
    rule_storage_write   => rule_writer_to_development_write,
    rule_storage_address => rule_writer_to_development_address,
    rule_storage_data    => rule_writer_to_development_data,

    decode_operation => decode_to_rule_writer_operation,
    decode_address   => decode_to_rule_writer_address,
    decode_data      => decode_to_rule_writer_data,

    run => run,

    clock => clock
  );

  development : entity work.development
  generic map (
    matrix_width             => matrix_width,
    matrix_height            => matrix_height,
    matrix_depth             => matrix_depth,
    matrix_wrap              => matrix_wrap,
    cell_type_bits           => cell_type_bits,
    cell_state_bits          => cell_state_bits,
    rule_amount              => rule_amount,
    rules_tested_in_parallel => rules_tested_in_parallel
  )
  port map (
    buffer_a_address_z    => development_to_mux_a_address_z,
    buffer_a_address_y    => development_to_mux_a_address_y,
    buffer_a_types_write  => development_to_mux_a_types_write,
    buffer_a_types_in     => development_from_mux_a_types,
    buffer_a_types_out    => development_to_mux_a_types,
    buffer_a_states_write => development_to_mux_a_states_write,
    buffer_a_states_in    => development_from_mux_a_states,
    buffer_a_states_out   => development_to_mux_a_states,

    buffer_b_address_z    => development_to_mux_b_address_z,
    buffer_b_address_y    => development_to_mux_b_address_y,
    buffer_b_types_write  => development_to_mux_b_types_write,
    buffer_b_types_in     => development_from_mux_b_types,
    buffer_b_types_out    => development_to_mux_b_types,
    buffer_b_states_write => development_to_mux_b_states_write,
    buffer_b_states_in    => development_from_mux_b_states,
    buffer_b_states_out   => development_to_mux_b_states,

    rule_storage_write   => rule_writer_to_development_write,
    rule_storage_address => rule_writer_to_development_address,
    rule_storage_data    => rule_writer_to_development_data,

    rule_vector_reader_data  => rule_vector_reader_from_development_data,
    rule_vector_reader_count => rule_vector_reader_from_development_count,
    rule_vector_reader_read  => rule_vector_reader_to_development_read,
    rule_vector_buffer_reset => decode_to_buffers_reset,

    rule_numbers_reader_address_z => rule_numbers_reader_to_development_address_z,
    rule_numbers_reader_address_y => rule_numbers_reader_to_development_address_y,
    rule_numbers_reader_data      => rule_numbers_reader_from_development_data,

    decode_operation    => decode_to_development_operation,
    decode_rules_active => decode_to_development_rules_active,

    run  => run,
    done => done_development,

    clock => clock
  );

  rule_vector_reader : entity work.rule_vector_reader
  generic map (
    rule_amount              => rule_amount,
    rule_vector_amount       => rule_vector_amount,
    send_buffer_address_bits => tx_buffer_address_bits
  )
  port map (
    vector_buffer_data  => rule_vector_reader_from_development_data,
    vector_buffer_count => rule_vector_reader_from_development_count,
    vector_buffer_read  => rule_vector_reader_to_development_read,

    send_buffer_data  => rule_vector_reader_to_send_mux_data,
    send_buffer_count => rule_vector_reader_from_send_mux_count,
    send_buffer_write => rule_vector_reader_to_send_mux_write,

    decode_operation => decode_to_rule_vector_reader_operation,
    decode_count     => decode_to_rule_vector_reader_count,

    run  => run,
    done => done_rule_vector_reader,

    clock => clock
  );

  rule_numbers_reader : entity work.rule_numbers_reader
  generic map (
    matrix_width             => matrix_width,
    matrix_height            => matrix_height,
    matrix_depth             => matrix_depth,
    rule_amount              => rule_amount,
    send_buffer_address_bits => tx_buffer_address_bits
  )
  port map (
    buffer_address_z => rule_numbers_reader_to_development_address_z,
    buffer_address_y => rule_numbers_reader_to_development_address_y,
    buffer_data      => rule_numbers_reader_from_development_data,

    send_buffer_data  => rule_numbers_reader_to_send_mux_data,
    send_buffer_count => rule_numbers_reader_from_send_mux_count,
    send_buffer_write => rule_numbers_reader_to_send_mux_write,

    decode_operation => decode_to_rule_numbers_reader_operation,

    run  => run,
    done => done_rule_numbers_reader,

    clock => clock
  );

  fitness : entity work.fitness_dft -- Change this to swap fitness module
  generic map (
    -- General fitness interface
    live_count_buffer_size => live_count_buffer_size,
    live_count_buffer_bits => live_count_buffer_bits,
    fitness_buffer_size    => fitness_buffer_size
    -- Spesific features are defined in each fitness module
  )
  port map (
    live_count_buffer_read  => fitness_to_live_count_buffer_read,
    live_count_buffer_data  => fitness_from_live_count_buffer_data,
    live_count_buffer_count => fitness_from_live_count_buffer_count,

    fitness_buffer_write => fitness_to_buffer_write,
    fitness_buffer_data  => fitness_to_buffer_data,
    fitness_buffer_count => fitness_buffer_count,

    identifier    => fitness_identifier,
    words_per_run => fitness_words_per_run,
    parameters    => fitness_parameters,

    clock => clock
  );

  fitness_buffer : entity work.fifo
  generic map (
    address_bits => bits(fitness_buffer_size),
    data_bits    => 32
  )
  port map (
    data_in    => fitness_to_buffer_data,
    data_out   => fitness_sender_from_buffer_data,
    data_count => fitness_buffer_count,
    data_read  => fitness_sender_to_buffer_read,
    data_write => fitness_to_buffer_write,
    reset      => decode_to_buffers_reset,
    clock      => clock
  );

  fitness_sender : entity work.fitness_sender
  generic map (
    send_buffer_size    => send_buffer_size,
    fitness_buffer_size => fitness_buffer_size
  )
  port map (
    send_buffer_write => fitness_sender_to_send_mux_write,
    send_buffer_data  => fitness_sender_to_send_mux_data,
    send_buffer_count => fitness_sender_from_send_mux_count,

    fitness_buffer_read  => fitness_sender_to_buffer_read,
    fitness_buffer_data  => fitness_sender_from_buffer_data,
    fitness_buffer_count => fitness_buffer_count,

    fitness_words_per_run => fitness_words_per_run,

    decode_operation => decode_to_fitness_sender_operation,

    run  => run,
    done => done_fitness_sender,

    clock => clock
  );

end rtl;
